New crossbar with Ideal transistors and big resistance range of memristors
$.option post ingold=1
.options post=2
.options MTTHRESH
.protect
.include '65nm_bulk.pm'
.hdl 'rram.va'
.unprotect

.param SET_PULSE=10ns   $ SET pulse width
.param SET_START=5ns    $ SET operation delay
.param RESET_PULSE=10ns $ RESET pulse width
.param RESET_START='SET_START+5n+SET_PULSE' $ RESET operation delay
.param T_FINAL='RESET_START+RESET_PULSE+5n' $ Final simulation time
.param V_0 = 0
.param V_1 = '1/3'
.param V_2 = '2/3'
.param V_3 = 1
.param Rmax=3e6
.param Rmin=10e3
.param Rf=10000
.param R =1000
.param RE='R/(Rf*(1/Rmin - 1/Rmax))'
.param ReOverR = '1/(Rf*(1/Rmin - 1/Rmax))'
.param gap_max=1.6693n
.param gap_min=0.1005n
.param gap_0 = gap_max
.param gap_1 = 0.4008n 
.param gap_2 = 0.2116n
.param gap_3 = gap_min


X1  BL1  SL1  rram    gap_ini=gap_3  tstep=10ps  $ RRAM1

X2  BL2  SL1  rram    gap_ini=gap_2  tstep=10ps  $ RRAM2

X3  BL3  SL1  rram    gap_ini=gap_1  tstep=10ps  $ RRAM3

X4  BL4  SL1  rram    gap_ini=gap_0  tstep=10ps  $ RRAM4

Xref1 BL1  SLref  rram    gap_ini=gap_max   tstep=10ps  $ RRAM reference 1
Xref2 BL2  SLref  rram    gap_ini=gap_max   tstep=10ps  $ RRAM reference 2
Xref3 BL3  SLref  rram    gap_ini=gap_max   tstep=10ps  $ RRAM reference 3
Xref4 BL4  SLref  rram    gap_ini=gap_max   tstep=10ps  $ RRAM reference 4

hV      V_SL     0 V_SL1_SET  Rf
hVref   V_Ref   0 V_SLref    Rf

e1      Vo    0 V_SL   V_Ref   ReOverR


V_Bias       Bias  0   PWL 0n 0
V_BL1        BL1   Bias   PWL (time, vol1)
V_BL2        BL2   Bias   PWL (time, vol2)
V_BL3        BL3   Bias   PWL (time, vol3)
V_BL4        BL4   Bias   PWL (time, vol4)
V_expected   expected 0   PWL (time, vol_exp)
.DATA vector
time vol1 vol2 vol3 vol4 vol_exp
0n 0.3333333333333333 1.0 0.0 1.0 1.0
9.999n 0.3333333333333333 1.0 0.0 1.0 1.0
10n 0.0 0.3333333333333333 1.0 0.3333333333333333 0.5555555555555556
19.999n 0.0 0.3333333333333333 1.0 0.3333333333333333 0.5555555555555556
20n 0.0 0.3333333333333333 1.0 1.0 0.5555555555555556
29.999n 0.0 0.3333333333333333 1.0 1.0 0.5555555555555556
30n 0.0 1.0 0.6666666666666666 0.0 0.8888888888888888
39.999n 0.0 1.0 0.6666666666666666 0.0 0.8888888888888888
40n 0.6666666666666666 0.0 1.0 0.3333333333333333 1.0
49.999n 0.6666666666666666 0.0 1.0 0.3333333333333333 1.0
50n 0.0 0.6666666666666666 0.0 1.0 0.4444444444444444
59.999n 0.0 0.6666666666666666 0.0 1.0 0.4444444444444444
60n 1.0 0.3333333333333333 0.3333333333333333 0.0 1.3333333333333333
69.999n 1.0 0.3333333333333333 0.3333333333333333 0.0 1.3333333333333333
70n 1.0 0.0 0.3333333333333333 0.3333333333333333 1.1111111111111112
79.999n 1.0 0.0 0.3333333333333333 0.3333333333333333 1.1111111111111112
80n 0.6666666666666666 0.0 1.0 1.0 1.0
89.999n 0.6666666666666666 0.0 1.0 1.0 1.0
90n 0.6666666666666666 1.0 0.0 0.6666666666666666 1.3333333333333333
99.999n 0.6666666666666666 1.0 0.0 0.6666666666666666 1.3333333333333333
100n 0.0 0.0 0.0 0.6666666666666666 0.0
109.999n 0.0 0.0 0.0 0.6666666666666666 0.0
110n 0.3333333333333333 1.0 0.0 1.0 1.0
119.999n 0.3333333333333333 1.0 0.0 1.0 1.0
120n 0.3333333333333333 0.6666666666666666 0.3333333333333333 0.3333333333333333 0.8888888888888888
129.999n 0.3333333333333333 0.6666666666666666 0.3333333333333333 0.3333333333333333 0.8888888888888888
130n 1.0 0.0 0.3333333333333333 0.6666666666666666 1.1111111111111112
139.999n 1.0 0.0 0.3333333333333333 0.6666666666666666 1.1111111111111112
140n 0.6666666666666666 1.0 0.3333333333333333 0.0 1.4444444444444444
149.999n 0.6666666666666666 1.0 0.3333333333333333 0.0 1.4444444444444444
150n 1.0 1.0 0.3333333333333333 1.0 1.7777777777777777
159.999n 1.0 1.0 0.3333333333333333 1.0 1.7777777777777777
160n 0.3333333333333333 0.3333333333333333 0.3333333333333333 0.6666666666666666 0.6666666666666666
169.999n 0.3333333333333333 0.3333333333333333 0.3333333333333333 0.6666666666666666 0.6666666666666666
170n 0.6666666666666666 1.0 0.0 0.6666666666666666 1.3333333333333333
179.999n 0.6666666666666666 1.0 0.0 0.6666666666666666 1.3333333333333333
180n 1.0 0.3333333333333333 0.3333333333333333 0.3333333333333333 1.3333333333333333
189.999n 1.0 0.3333333333333333 0.3333333333333333 0.3333333333333333 1.3333333333333333
190n 0.3333333333333333 0.0 1.0 0.3333333333333333 0.6666666666666666
199.999n 0.3333333333333333 0.0 1.0 0.3333333333333333 0.6666666666666666
200n 0.3333333333333333 0.3333333333333333 1.0 0.0 0.8888888888888888
209.999n 0.3333333333333333 0.3333333333333333 1.0 0.0 0.8888888888888888
210n 0.0 1.0 0.6666666666666666 0.6666666666666666 0.8888888888888888
219.999n 0.0 1.0 0.6666666666666666 0.6666666666666666 0.8888888888888888
220n 0.6666666666666666 0.0 1.0 1.0 1.0
229.999n 0.6666666666666666 0.0 1.0 1.0 1.0
230n 1.0 1.0 1.0 0.0 2.0
239.999n 1.0 1.0 1.0 0.0 2.0
240n 0.6666666666666666 0.0 0.6666666666666666 0.0 0.8888888888888888
249.999n 0.6666666666666666 0.0 0.6666666666666666 0.0 0.8888888888888888
250n 0.3333333333333333 1.0 1.0 1.0 1.3333333333333333
259.999n 0.3333333333333333 1.0 1.0 1.0 1.3333333333333333
260n 0.6666666666666666 0.0 0.3333333333333333 0.3333333333333333 0.7777777777777778
269.999n 0.6666666666666666 0.0 0.3333333333333333 0.3333333333333333 0.7777777777777778
270n 0.3333333333333333 1.0 1.0 0.0 1.3333333333333333
279.999n 0.3333333333333333 1.0 1.0 0.0 1.3333333333333333
280n 0.0 0.3333333333333333 0.3333333333333333 0.3333333333333333 0.3333333333333333
289.999n 0.0 0.3333333333333333 0.3333333333333333 0.3333333333333333 0.3333333333333333
290n 0.6666666666666666 1.0 0.6666666666666666 0.6666666666666666 1.5555555555555556
299.999n 0.6666666666666666 1.0 0.6666666666666666 0.6666666666666666 1.5555555555555556
300n 1.0 0.6666666666666666 1.0 0.3333333333333333 1.7777777777777777
309.999n 1.0 0.6666666666666666 1.0 0.3333333333333333 1.7777777777777777
310n 1.0 0.0 1.0 0.3333333333333333 1.3333333333333333
319.999n 1.0 0.0 1.0 0.3333333333333333 1.3333333333333333
320n 0.0 0.0 1.0 1.0 0.3333333333333333
329.999n 0.0 0.0 1.0 1.0 0.3333333333333333
330n 0.0 0.0 0.0 0.3333333333333333 0.0
339.999n 0.0 0.0 0.0 0.3333333333333333 0.0
340n 1.0 1.0 0.0 0.0 1.6666666666666667
349.999n 1.0 1.0 0.0 0.0 1.6666666666666667
350n 1.0 1.0 1.0 0.6666666666666666 2.0
359.999n 1.0 1.0 1.0 0.6666666666666666 2.0
360n 0.0 0.3333333333333333 0.3333333333333333 1.0 0.3333333333333333
369.999n 0.0 0.3333333333333333 0.3333333333333333 1.0 0.3333333333333333
370n 0.6666666666666666 0.3333333333333333 0.0 1.0 0.8888888888888888
379.999n 0.6666666666666666 0.3333333333333333 0.0 1.0 0.8888888888888888
380n 0.3333333333333333 0.6666666666666666 0.6666666666666666 0.0 1.0
389.999n 0.3333333333333333 0.6666666666666666 0.6666666666666666 0.0 1.0
390n 0.0 1.0 0.0 0.0 0.6666666666666666
399.999n 0.0 1.0 0.0 0.0 0.6666666666666666
400n 0.0 0.3333333333333333 0.6666666666666666 0.6666666666666666 0.4444444444444444
409.999n 0.0 0.3333333333333333 0.6666666666666666 0.6666666666666666 0.4444444444444444
410n 0.0 1.0 0.0 1.0 0.6666666666666666
419.999n 0.0 1.0 0.0 1.0 0.6666666666666666
420n 0.3333333333333333 1.0 0.0 1.0 1.0
429.999n 0.3333333333333333 1.0 0.0 1.0 1.0
430n 0.0 0.3333333333333333 1.0 0.3333333333333333 0.5555555555555556
439.999n 0.0 0.3333333333333333 1.0 0.3333333333333333 0.5555555555555556
440n 1.0 0.3333333333333333 1.0 1.0 1.5555555555555556
449.999n 1.0 0.3333333333333333 1.0 1.0 1.5555555555555556
450n 0.6666666666666666 0.6666666666666666 0.6666666666666666 0.0 1.3333333333333333
459.999n 0.6666666666666666 0.6666666666666666 0.6666666666666666 0.0 1.3333333333333333
460n 0.6666666666666666 0.0 0.0 0.0 0.6666666666666666
469.999n 0.6666666666666666 0.0 0.0 0.0 0.6666666666666666
470n 0.6666666666666666 0.6666666666666666 0.0 0.0 1.1111111111111112
479.999n 0.6666666666666666 0.6666666666666666 0.0 0.0 1.1111111111111112
480n 0.0 1.0 1.0 1.0 1.0
489.999n 0.0 1.0 1.0 1.0 1.0
490n 0.0 0.6666666666666666 1.0 1.0 0.7777777777777778
499.999n 0.0 0.6666666666666666 1.0 1.0 0.7777777777777778
500n 1.0 1.0 0.3333333333333333 0.0 1.7777777777777777
509.999n 1.0 1.0 0.3333333333333333 0.0 1.7777777777777777
510n 0.0 0.3333333333333333 1.0 0.3333333333333333 0.5555555555555556
519.999n 0.0 0.3333333333333333 1.0 0.3333333333333333 0.5555555555555556
520n 1.0 0.3333333333333333 0.3333333333333333 0.3333333333333333 1.3333333333333333
529.999n 1.0 0.3333333333333333 0.3333333333333333 0.3333333333333333 1.3333333333333333
530n 0.0 0.3333333333333333 0.0 0.3333333333333333 0.2222222222222222
539.999n 0.0 0.3333333333333333 0.0 0.3333333333333333 0.2222222222222222
540n 1.0 0.3333333333333333 1.0 1.0 1.5555555555555556
549.999n 1.0 0.3333333333333333 1.0 1.0 1.5555555555555556
550n 0.6666666666666666 1.0 0.0 0.6666666666666666 1.3333333333333333
559.999n 0.6666666666666666 1.0 0.0 0.6666666666666666 1.3333333333333333
560n 1.0 0.3333333333333333 0.6666666666666666 0.6666666666666666 1.4444444444444444
569.999n 1.0 0.3333333333333333 0.6666666666666666 0.6666666666666666 1.4444444444444444
570n 0.3333333333333333 0.0 0.0 0.6666666666666666 0.3333333333333333
579.999n 0.3333333333333333 0.0 0.0 0.6666666666666666 0.3333333333333333
580n 1.0 0.0 0.6666666666666666 1.0 1.2222222222222223
589.999n 1.0 0.0 0.6666666666666666 1.0 1.2222222222222223
590n 0.0 0.0 0.3333333333333333 0.3333333333333333 0.1111111111111111
599.999n 0.0 0.0 0.3333333333333333 0.3333333333333333 0.1111111111111111
600n 0.3333333333333333 0.0 1.0 0.3333333333333333 0.6666666666666666
609.999n 0.3333333333333333 0.0 1.0 0.3333333333333333 0.6666666666666666
610n 0.3333333333333333 0.6666666666666666 0.3333333333333333 1.0 0.8888888888888888
619.999n 0.3333333333333333 0.6666666666666666 0.3333333333333333 1.0 0.8888888888888888
620n 0.0 0.3333333333333333 1.0 0.0 0.5555555555555556
629.999n 0.0 0.3333333333333333 1.0 0.0 0.5555555555555556
630n 0.6666666666666666 0.6666666666666666 0.3333333333333333 1.0 1.2222222222222223
639.999n 0.6666666666666666 0.6666666666666666 0.3333333333333333 1.0 1.2222222222222223
640n 0.0 0.3333333333333333 0.0 1.0 0.2222222222222222
649.999n 0.0 0.3333333333333333 0.0 1.0 0.2222222222222222
650n 0.6666666666666666 0.6666666666666666 0.3333333333333333 0.3333333333333333 1.2222222222222223
659.999n 0.6666666666666666 0.6666666666666666 0.3333333333333333 0.3333333333333333 1.2222222222222223
660n 0.3333333333333333 0.3333333333333333 1.0 0.0 0.8888888888888888
669.999n 0.3333333333333333 0.3333333333333333 1.0 0.0 0.8888888888888888
670n 0.6666666666666666 0.0 1.0 1.0 1.0
679.999n 0.6666666666666666 0.0 1.0 1.0 1.0
680n 0.6666666666666666 0.6666666666666666 0.6666666666666666 1.0 1.3333333333333333
689.999n 0.6666666666666666 0.6666666666666666 0.6666666666666666 1.0 1.3333333333333333
690n 0.3333333333333333 0.6666666666666666 0.0 1.0 0.7777777777777778
699.999n 0.3333333333333333 0.6666666666666666 0.0 1.0 0.7777777777777778
700n 0.6666666666666666 1.0 1.0 0.0 1.6666666666666667
709.999n 0.6666666666666666 1.0 1.0 0.0 1.6666666666666667
710n 0.6666666666666666 0.6666666666666666 0.3333333333333333 0.6666666666666666 1.2222222222222223
719.999n 0.6666666666666666 0.6666666666666666 0.3333333333333333 0.6666666666666666 1.2222222222222223
720n 0.0 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.5555555555555556
729.999n 0.0 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.5555555555555556
730n 0.6666666666666666 0.3333333333333333 0.3333333333333333 0.0 1.0
739.999n 0.6666666666666666 0.3333333333333333 0.3333333333333333 0.0 1.0
740n 0.0 0.3333333333333333 1.0 0.0 0.5555555555555556
749.999n 0.0 0.3333333333333333 1.0 0.0 0.5555555555555556
750n 0.3333333333333333 0.6666666666666666 0.0 1.0 0.7777777777777778
759.999n 0.3333333333333333 0.6666666666666666 0.0 1.0 0.7777777777777778
760n 0.3333333333333333 1.0 1.0 0.0 1.3333333333333333
769.999n 0.3333333333333333 1.0 1.0 0.0 1.3333333333333333
770n 0.6666666666666666 0.0 1.0 1.0 1.0
779.999n 0.6666666666666666 0.0 1.0 1.0 1.0
780n 0.0 0.6666666666666666 0.6666666666666666 0.6666666666666666 0.6666666666666666
789.999n 0.0 0.6666666666666666 0.6666666666666666 0.6666666666666666 0.6666666666666666
790n 0.3333333333333333 0.0 0.6666666666666666 0.3333333333333333 0.5555555555555556
799.999n 0.3333333333333333 0.0 0.6666666666666666 0.3333333333333333 0.5555555555555556
800n 0.3333333333333333 1.0 0.6666666666666666 0.3333333333333333 1.2222222222222223
809.999n 0.3333333333333333 1.0 0.6666666666666666 0.3333333333333333 1.2222222222222223
810n 0.3333333333333333 0.6666666666666666 1.0 0.0 1.1111111111111112
819.999n 0.3333333333333333 0.6666666666666666 1.0 0.0 1.1111111111111112
820n 0.6666666666666666 0.0 0.0 0.0 0.6666666666666666
829.999n 0.6666666666666666 0.0 0.0 0.0 0.6666666666666666
830n 0.3333333333333333 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.8888888888888888
839.999n 0.3333333333333333 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.8888888888888888
840n 0.0 1.0 1.0 0.6666666666666666 1.0
849.999n 0.0 1.0 1.0 0.6666666666666666 1.0
850n 0.0 0.3333333333333333 0.6666666666666666 0.0 0.4444444444444444
859.999n 0.0 0.3333333333333333 0.6666666666666666 0.0 0.4444444444444444
860n 1.0 0.3333333333333333 0.0 1.0 1.2222222222222223
869.999n 1.0 0.3333333333333333 0.0 1.0 1.2222222222222223
870n 0.0 0.3333333333333333 0.6666666666666666 1.0 0.4444444444444444
879.999n 0.0 0.3333333333333333 0.6666666666666666 1.0 0.4444444444444444
880n 0.6666666666666666 0.3333333333333333 0.3333333333333333 0.6666666666666666 1.0
889.999n 0.6666666666666666 0.3333333333333333 0.3333333333333333 0.6666666666666666 1.0
890n 0.6666666666666666 0.6666666666666666 1.0 0.6666666666666666 1.4444444444444444
899.999n 0.6666666666666666 0.6666666666666666 1.0 0.6666666666666666 1.4444444444444444
900n 0.0 0.6666666666666666 0.3333333333333333 0.0 0.5555555555555556
909.999n 0.0 0.6666666666666666 0.3333333333333333 0.0 0.5555555555555556
910n 0.0 1.0 1.0 0.6666666666666666 1.0
919.999n 0.0 1.0 1.0 0.6666666666666666 1.0
920n 1.0 1.0 0.0 0.0 1.6666666666666667
929.999n 1.0 1.0 0.0 0.0 1.6666666666666667
930n 0.0 1.0 0.6666666666666666 1.0 0.8888888888888888
939.999n 0.0 1.0 0.6666666666666666 1.0 0.8888888888888888
940n 0.3333333333333333 0.0 0.0 1.0 0.3333333333333333
949.999n 0.3333333333333333 0.0 0.0 1.0 0.3333333333333333
950n 0.3333333333333333 0.0 0.6666666666666666 0.0 0.5555555555555556
959.999n 0.3333333333333333 0.0 0.6666666666666666 0.0 0.5555555555555556
960n 0.0 0.0 1.0 0.0 0.3333333333333333
969.999n 0.0 0.0 1.0 0.0 0.3333333333333333
970n 0.0 0.6666666666666666 0.0 0.3333333333333333 0.4444444444444444
979.999n 0.0 0.6666666666666666 0.0 0.3333333333333333 0.4444444444444444
980n 0.6666666666666666 0.0 0.3333333333333333 0.6666666666666666 0.7777777777777778
989.999n 0.6666666666666666 0.0 0.3333333333333333 0.6666666666666666 0.7777777777777778
990n 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.6666666666666666 1.1111111111111112
999.999n 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.6666666666666666 1.1111111111111112
1000n 0.0 0.3333333333333333 1.0 1.0 0.5555555555555556
1009.999n 0.0 0.3333333333333333 1.0 1.0 0.5555555555555556
1010n 0.6666666666666666 0.0 0.6666666666666666 0.6666666666666666 0.8888888888888888
1019.999n 0.6666666666666666 0.0 0.6666666666666666 0.6666666666666666 0.8888888888888888
1020n 0.0 0.6666666666666666 0.0 0.3333333333333333 0.4444444444444444
1029.999n 0.0 0.6666666666666666 0.0 0.3333333333333333 0.4444444444444444
1030n 0.3333333333333333 0.0 1.0 0.0 0.6666666666666666
1039.999n 0.3333333333333333 0.0 1.0 0.0 0.6666666666666666
1040n 0.0 1.0 0.6666666666666666 0.6666666666666666 0.8888888888888888
1049.999n 0.0 1.0 0.6666666666666666 0.6666666666666666 0.8888888888888888
1050n 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.6666666666666666 1.1111111111111112
1059.999n 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.6666666666666666 1.1111111111111112
1060n 0.6666666666666666 1.0 1.0 0.6666666666666666 1.6666666666666667
1069.999n 0.6666666666666666 1.0 1.0 0.6666666666666666 1.6666666666666667
1070n 1.0 0.0 1.0 0.6666666666666666 1.3333333333333333
1079.999n 1.0 0.0 1.0 0.6666666666666666 1.3333333333333333
1080n 1.0 1.0 0.6666666666666666 1.0 1.8888888888888888
1089.999n 1.0 1.0 0.6666666666666666 1.0 1.8888888888888888
1090n 0.6666666666666666 1.0 1.0 0.3333333333333333 1.6666666666666667
1099.999n 0.6666666666666666 1.0 1.0 0.3333333333333333 1.6666666666666667
1100n 0.3333333333333333 0.0 0.6666666666666666 0.0 0.5555555555555556
1109.999n 0.3333333333333333 0.0 0.6666666666666666 0.0 0.5555555555555556
1110n 1.0 1.0 0.3333333333333333 0.6666666666666666 1.7777777777777777
1119.999n 1.0 1.0 0.3333333333333333 0.6666666666666666 1.7777777777777777
1120n 1.0 0.6666666666666666 1.0 0.0 1.7777777777777777
1129.999n 1.0 0.6666666666666666 1.0 0.0 1.7777777777777777
1130n 0.0 1.0 0.3333333333333333 1.0 0.7777777777777778
1139.999n 0.0 1.0 0.3333333333333333 1.0 0.7777777777777778
1140n 1.0 1.0 0.3333333333333333 0.6666666666666666 1.7777777777777777
1149.999n 1.0 1.0 0.3333333333333333 0.6666666666666666 1.7777777777777777
1150n 0.0 1.0 1.0 0.0 1.0
1159.999n 0.0 1.0 1.0 0.0 1.0
1160n 0.3333333333333333 0.3333333333333333 0.6666666666666666 0.0 0.7777777777777778
1169.999n 0.3333333333333333 0.3333333333333333 0.6666666666666666 0.0 0.7777777777777778
1170n 0.0 1.0 1.0 0.0 1.0
1179.999n 0.0 1.0 1.0 0.0 1.0
1180n 1.0 0.0 1.0 0.3333333333333333 1.3333333333333333
1189.999n 1.0 0.0 1.0 0.3333333333333333 1.3333333333333333
1190n 1.0 0.0 0.6666666666666666 0.3333333333333333 1.2222222222222223
1199.999n 1.0 0.0 0.6666666666666666 0.3333333333333333 1.2222222222222223
1200n 1.0 0.6666666666666666 0.0 0.0 1.4444444444444444
1209.999n 1.0 0.6666666666666666 0.0 0.0 1.4444444444444444
1210n 0.6666666666666666 1.0 0.0 0.3333333333333333 1.3333333333333333
1219.999n 0.6666666666666666 1.0 0.0 0.3333333333333333 1.3333333333333333
1220n 0.6666666666666666 0.3333333333333333 0.0 0.0 0.8888888888888888
1229.999n 0.6666666666666666 0.3333333333333333 0.0 0.0 0.8888888888888888
1230n 0.0 0.3333333333333333 0.3333333333333333 0.6666666666666666 0.3333333333333333
1239.999n 0.0 0.3333333333333333 0.3333333333333333 0.6666666666666666 0.3333333333333333
1240n 0.0 0.3333333333333333 0.3333333333333333 0.6666666666666666 0.3333333333333333
1249.999n 0.0 0.3333333333333333 0.3333333333333333 0.6666666666666666 0.3333333333333333
1250n 0.6666666666666666 1.0 0.0 1.0 1.3333333333333333
1259.999n 0.6666666666666666 1.0 0.0 1.0 1.3333333333333333
1260n 0.6666666666666666 0.6666666666666666 0.3333333333333333 0.0 1.2222222222222223
1269.999n 0.6666666666666666 0.6666666666666666 0.3333333333333333 0.0 1.2222222222222223
1270n 1.0 0.3333333333333333 1.0 0.6666666666666666 1.5555555555555556
1279.999n 1.0 0.3333333333333333 1.0 0.6666666666666666 1.5555555555555556
1280n 0.6666666666666666 1.0 1.0 0.0 1.6666666666666667
1289.999n 0.6666666666666666 1.0 1.0 0.0 1.6666666666666667
1290n 0.3333333333333333 0.0 0.3333333333333333 0.6666666666666666 0.4444444444444444
1299.999n 0.3333333333333333 0.0 0.3333333333333333 0.6666666666666666 0.4444444444444444
1300n 1.0 0.3333333333333333 0.0 0.0 1.2222222222222223
1309.999n 1.0 0.3333333333333333 0.0 0.0 1.2222222222222223
1310n 1.0 0.0 1.0 0.3333333333333333 1.3333333333333333
1319.999n 1.0 0.0 1.0 0.3333333333333333 1.3333333333333333
1320n 0.0 1.0 0.3333333333333333 0.0 0.7777777777777778
1329.999n 0.0 1.0 0.3333333333333333 0.0 0.7777777777777778
1330n 1.0 1.0 0.0 0.6666666666666666 1.6666666666666667
1339.999n 1.0 1.0 0.0 0.6666666666666666 1.6666666666666667
1340n 0.3333333333333333 0.6666666666666666 1.0 1.0 1.1111111111111112
1349.999n 0.3333333333333333 0.6666666666666666 1.0 1.0 1.1111111111111112
1350n 0.6666666666666666 0.0 0.0 1.0 0.6666666666666666
1359.999n 0.6666666666666666 0.0 0.0 1.0 0.6666666666666666
1360n 0.0 0.6666666666666666 0.0 0.0 0.4444444444444444
1369.999n 0.0 0.6666666666666666 0.0 0.0 0.4444444444444444
1370n 1.0 0.6666666666666666 0.3333333333333333 1.0 1.5555555555555556
1379.999n 1.0 0.6666666666666666 0.3333333333333333 1.0 1.5555555555555556
1380n 0.0 0.0 1.0 1.0 0.3333333333333333
1389.999n 0.0 0.0 1.0 1.0 0.3333333333333333
1390n 0.3333333333333333 0.3333333333333333 0.3333333333333333 0.6666666666666666 0.6666666666666666
1399.999n 0.3333333333333333 0.3333333333333333 0.3333333333333333 0.6666666666666666 0.6666666666666666
1400n 0.6666666666666666 0.6666666666666666 0.3333333333333333 0.0 1.2222222222222223
1409.999n 0.6666666666666666 0.6666666666666666 0.3333333333333333 0.0 1.2222222222222223
1410n 0.6666666666666666 0.3333333333333333 1.0 0.3333333333333333 1.2222222222222223
1419.999n 0.6666666666666666 0.3333333333333333 1.0 0.3333333333333333 1.2222222222222223
1420n 1.0 0.3333333333333333 1.0 0.0 1.5555555555555556
1429.999n 1.0 0.3333333333333333 1.0 0.0 1.5555555555555556
1430n 0.3333333333333333 0.0 1.0 0.6666666666666666 0.6666666666666666
1439.999n 0.3333333333333333 0.0 1.0 0.6666666666666666 0.6666666666666666
1440n 0.3333333333333333 0.0 1.0 0.0 0.6666666666666666
1449.999n 0.3333333333333333 0.0 1.0 0.0 0.6666666666666666
1450n 0.3333333333333333 0.6666666666666666 0.0 0.3333333333333333 0.7777777777777778
1459.999n 0.3333333333333333 0.6666666666666666 0.0 0.3333333333333333 0.7777777777777778
1460n 0.0 0.3333333333333333 0.3333333333333333 0.0 0.3333333333333333
1469.999n 0.0 0.3333333333333333 0.3333333333333333 0.0 0.3333333333333333
1470n 0.6666666666666666 0.0 0.6666666666666666 0.3333333333333333 0.8888888888888888
1479.999n 0.6666666666666666 0.0 0.6666666666666666 0.3333333333333333 0.8888888888888888
1480n 0.6666666666666666 0.6666666666666666 1.0 0.6666666666666666 1.4444444444444444
1489.999n 0.6666666666666666 0.6666666666666666 1.0 0.6666666666666666 1.4444444444444444
1490n 0.6666666666666666 1.0 0.6666666666666666 0.6666666666666666 1.5555555555555556
1499.999n 0.6666666666666666 1.0 0.6666666666666666 0.6666666666666666 1.5555555555555556
1500n 0.0 0.6666666666666666 0.0 0.0 0.4444444444444444
1509.999n 0.0 0.6666666666666666 0.0 0.0 0.4444444444444444
1510n 1.0 0.0 0.0 0.3333333333333333 1.0
1519.999n 1.0 0.0 0.0 0.3333333333333333 1.0
1520n 0.6666666666666666 0.0 0.3333333333333333 0.0 0.7777777777777778
1529.999n 0.6666666666666666 0.0 0.3333333333333333 0.0 0.7777777777777778
1530n 0.0 0.3333333333333333 0.3333333333333333 0.3333333333333333 0.3333333333333333
1539.999n 0.0 0.3333333333333333 0.3333333333333333 0.3333333333333333 0.3333333333333333
1540n 0.3333333333333333 0.0 0.6666666666666666 0.0 0.5555555555555556
1549.999n 0.3333333333333333 0.0 0.6666666666666666 0.0 0.5555555555555556
1550n 0.3333333333333333 1.0 1.0 1.0 1.3333333333333333
1559.999n 0.3333333333333333 1.0 1.0 1.0 1.3333333333333333
1560n 0.6666666666666666 0.3333333333333333 0.0 0.3333333333333333 0.8888888888888888
1569.999n 0.6666666666666666 0.3333333333333333 0.0 0.3333333333333333 0.8888888888888888
1570n 1.0 0.3333333333333333 0.0 1.0 1.2222222222222223
1579.999n 1.0 0.3333333333333333 0.0 1.0 1.2222222222222223
1580n 0.3333333333333333 0.6666666666666666 0.0 1.0 0.7777777777777778
1589.999n 0.3333333333333333 0.6666666666666666 0.0 1.0 0.7777777777777778
1590n 0.0 0.0 1.0 1.0 0.3333333333333333
1599.999n 0.0 0.0 1.0 1.0 0.3333333333333333
1600n 0.6666666666666666 0.3333333333333333 1.0 0.6666666666666666 1.2222222222222223
1609.999n 0.6666666666666666 0.3333333333333333 1.0 0.6666666666666666 1.2222222222222223
1610n 0.6666666666666666 1.0 0.6666666666666666 0.0 1.5555555555555556
1619.999n 0.6666666666666666 1.0 0.6666666666666666 0.0 1.5555555555555556
1620n 0.3333333333333333 1.0 0.0 0.6666666666666666 1.0
1629.999n 0.3333333333333333 1.0 0.0 0.6666666666666666 1.0
1630n 0.6666666666666666 1.0 0.3333333333333333 0.6666666666666666 1.4444444444444444
1639.999n 0.6666666666666666 1.0 0.3333333333333333 0.6666666666666666 1.4444444444444444
1640n 0.3333333333333333 0.0 0.6666666666666666 0.6666666666666666 0.5555555555555556
1649.999n 0.3333333333333333 0.0 0.6666666666666666 0.6666666666666666 0.5555555555555556
1650n 0.3333333333333333 0.3333333333333333 0.3333333333333333 0.3333333333333333 0.6666666666666666
1659.999n 0.3333333333333333 0.3333333333333333 0.3333333333333333 0.3333333333333333 0.6666666666666666
1660n 0.3333333333333333 0.0 1.0 0.6666666666666666 0.6666666666666666
1669.999n 0.3333333333333333 0.0 1.0 0.6666666666666666 0.6666666666666666
1670n 0.0 0.3333333333333333 0.0 0.6666666666666666 0.2222222222222222
1679.999n 0.0 0.3333333333333333 0.0 0.6666666666666666 0.2222222222222222
1680n 0.6666666666666666 0.0 0.6666666666666666 1.0 0.8888888888888888
1689.999n 0.6666666666666666 0.0 0.6666666666666666 1.0 0.8888888888888888
1690n 0.6666666666666666 0.3333333333333333 0.3333333333333333 1.0 1.0
1699.999n 0.6666666666666666 0.3333333333333333 0.3333333333333333 1.0 1.0
1700n 0.0 0.6666666666666666 0.3333333333333333 0.0 0.5555555555555556
1709.999n 0.0 0.6666666666666666 0.3333333333333333 0.0 0.5555555555555556
1710n 0.0 0.0 0.6666666666666666 0.0 0.2222222222222222
1719.999n 0.0 0.0 0.6666666666666666 0.0 0.2222222222222222
1720n 0.0 0.0 0.6666666666666666 1.0 0.2222222222222222
1729.999n 0.0 0.0 0.6666666666666666 1.0 0.2222222222222222
1730n 0.6666666666666666 1.0 0.6666666666666666 0.0 1.5555555555555556
1739.999n 0.6666666666666666 1.0 0.6666666666666666 0.0 1.5555555555555556
1740n 0.0 1.0 1.0 0.0 1.0
1749.999n 0.0 1.0 1.0 0.0 1.0
1750n 0.3333333333333333 1.0 0.6666666666666666 0.6666666666666666 1.2222222222222223
1759.999n 0.3333333333333333 1.0 0.6666666666666666 0.6666666666666666 1.2222222222222223
1760n 1.0 0.0 0.6666666666666666 1.0 1.2222222222222223
1769.999n 1.0 0.0 0.6666666666666666 1.0 1.2222222222222223
1770n 0.0 0.6666666666666666 0.0 0.6666666666666666 0.4444444444444444
1779.999n 0.0 0.6666666666666666 0.0 0.6666666666666666 0.4444444444444444
1780n 0.6666666666666666 0.6666666666666666 0.3333333333333333 0.0 1.2222222222222223
1789.999n 0.6666666666666666 0.6666666666666666 0.3333333333333333 0.0 1.2222222222222223
1790n 0.6666666666666666 1.0 1.0 0.6666666666666666 1.6666666666666667
1799.999n 0.6666666666666666 1.0 1.0 0.6666666666666666 1.6666666666666667
1800n 0.6666666666666666 0.6666666666666666 0.6666666666666666 0.3333333333333333 1.3333333333333333
1809.999n 0.6666666666666666 0.6666666666666666 0.6666666666666666 0.3333333333333333 1.3333333333333333
1810n 1.0 1.0 0.6666666666666666 0.3333333333333333 1.8888888888888888
1819.999n 1.0 1.0 0.6666666666666666 0.3333333333333333 1.8888888888888888
1820n 0.3333333333333333 0.6666666666666666 1.0 0.3333333333333333 1.1111111111111112
1829.999n 0.3333333333333333 0.6666666666666666 1.0 0.3333333333333333 1.1111111111111112
1830n 0.3333333333333333 0.3333333333333333 0.6666666666666666 0.3333333333333333 0.7777777777777778
1839.999n 0.3333333333333333 0.3333333333333333 0.6666666666666666 0.3333333333333333 0.7777777777777778
1840n 0.6666666666666666 1.0 0.6666666666666666 0.6666666666666666 1.5555555555555556
1849.999n 0.6666666666666666 1.0 0.6666666666666666 0.6666666666666666 1.5555555555555556
1850n 0.6666666666666666 0.3333333333333333 0.0 1.0 0.8888888888888888
1859.999n 0.6666666666666666 0.3333333333333333 0.0 1.0 0.8888888888888888
1860n 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.6666666666666666 1.1111111111111112
1869.999n 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.6666666666666666 1.1111111111111112
1870n 1.0 0.3333333333333333 0.0 0.3333333333333333 1.2222222222222223
1879.999n 1.0 0.3333333333333333 0.0 0.3333333333333333 1.2222222222222223
1880n 0.0 1.0 0.0 0.0 0.6666666666666666
1889.999n 0.0 1.0 0.0 0.0 0.6666666666666666
1890n 0.3333333333333333 0.3333333333333333 0.3333333333333333 0.0 0.6666666666666666
1899.999n 0.3333333333333333 0.3333333333333333 0.3333333333333333 0.0 0.6666666666666666
1900n 0.3333333333333333 1.0 1.0 0.6666666666666666 1.3333333333333333
1909.999n 0.3333333333333333 1.0 1.0 0.6666666666666666 1.3333333333333333
1910n 0.6666666666666666 0.0 1.0 0.6666666666666666 1.0
1919.999n 0.6666666666666666 0.0 1.0 0.6666666666666666 1.0
1920n 1.0 0.6666666666666666 0.6666666666666666 0.0 1.6666666666666667
1929.999n 1.0 0.6666666666666666 0.6666666666666666 0.0 1.6666666666666667
1930n 0.0 0.0 0.0 0.0 0.0
1939.999n 0.0 0.0 0.0 0.0 0.0
1940n 0.0 0.3333333333333333 0.6666666666666666 0.0 0.4444444444444444
1949.999n 0.0 0.3333333333333333 0.6666666666666666 0.0 0.4444444444444444
1950n 1.0 1.0 0.0 0.0 1.6666666666666667
1959.999n 1.0 1.0 0.0 0.0 1.6666666666666667
1960n 0.3333333333333333 0.0 0.6666666666666666 0.3333333333333333 0.5555555555555556
1969.999n 0.3333333333333333 0.0 0.6666666666666666 0.3333333333333333 0.5555555555555556
1970n 0.3333333333333333 0.6666666666666666 0.3333333333333333 0.0 0.8888888888888888
1979.999n 0.3333333333333333 0.6666666666666666 0.3333333333333333 0.0 0.8888888888888888
1980n 1.0 0.3333333333333333 1.0 0.6666666666666666 1.5555555555555556
1989.999n 1.0 0.3333333333333333 1.0 0.6666666666666666 1.5555555555555556
1990n 1.0 0.6666666666666666 0.6666666666666666 0.3333333333333333 1.6666666666666667
1999.999n 1.0 0.6666666666666666 0.6666666666666666 0.3333333333333333 1.6666666666666667
2000n 1.0 0.0 1.0 1.0 1.3333333333333333
2009.999n 1.0 0.0 1.0 1.0 1.3333333333333333
2010n 1.0 0.3333333333333333 0.6666666666666666 0.6666666666666666 1.4444444444444444
2019.999n 1.0 0.3333333333333333 0.6666666666666666 0.6666666666666666 1.4444444444444444
2020n 0.6666666666666666 0.0 0.3333333333333333 0.3333333333333333 0.7777777777777778
2029.999n 0.6666666666666666 0.0 0.3333333333333333 0.3333333333333333 0.7777777777777778
2030n 0.6666666666666666 0.0 1.0 0.0 1.0
2039.999n 0.6666666666666666 0.0 1.0 0.0 1.0
2040n 0.0 1.0 0.3333333333333333 0.0 0.7777777777777778
2049.999n 0.0 1.0 0.3333333333333333 0.0 0.7777777777777778
2050n 0.3333333333333333 0.3333333333333333 0.3333333333333333 1.0 0.6666666666666666
2059.999n 0.3333333333333333 0.3333333333333333 0.3333333333333333 1.0 0.6666666666666666
2060n 0.0 1.0 1.0 0.6666666666666666 1.0
2069.999n 0.0 1.0 1.0 0.6666666666666666 1.0
2070n 0.6666666666666666 0.0 1.0 1.0 1.0
2079.999n 0.6666666666666666 0.0 1.0 1.0 1.0
2080n 0.6666666666666666 0.3333333333333333 0.6666666666666666 1.0 1.1111111111111112
2089.999n 0.6666666666666666 0.3333333333333333 0.6666666666666666 1.0 1.1111111111111112
2090n 0.0 1.0 0.6666666666666666 0.3333333333333333 0.8888888888888888
2099.999n 0.0 1.0 0.6666666666666666 0.3333333333333333 0.8888888888888888
2100n 0.6666666666666666 0.6666666666666666 0.3333333333333333 0.3333333333333333 1.2222222222222223
2109.999n 0.6666666666666666 0.6666666666666666 0.3333333333333333 0.3333333333333333 1.2222222222222223
2110n 0.0 0.3333333333333333 0.6666666666666666 1.0 0.4444444444444444
2119.999n 0.0 0.3333333333333333 0.6666666666666666 1.0 0.4444444444444444
2120n 0.0 0.3333333333333333 1.0 0.0 0.5555555555555556
2129.999n 0.0 0.3333333333333333 1.0 0.0 0.5555555555555556
2130n 0.6666666666666666 0.6666666666666666 0.0 0.3333333333333333 1.1111111111111112
2139.999n 0.6666666666666666 0.6666666666666666 0.0 0.3333333333333333 1.1111111111111112
2140n 0.0 1.0 0.3333333333333333 0.0 0.7777777777777778
2149.999n 0.0 1.0 0.3333333333333333 0.0 0.7777777777777778
2150n 0.0 1.0 0.0 0.6666666666666666 0.6666666666666666
2159.999n 0.0 1.0 0.0 0.6666666666666666 0.6666666666666666
2160n 0.3333333333333333 1.0 0.3333333333333333 1.0 1.1111111111111112
2169.999n 0.3333333333333333 1.0 0.3333333333333333 1.0 1.1111111111111112
2170n 0.0 1.0 0.6666666666666666 1.0 0.8888888888888888
2179.999n 0.0 1.0 0.6666666666666666 1.0 0.8888888888888888
2180n 0.0 0.3333333333333333 0.6666666666666666 0.3333333333333333 0.4444444444444444
2189.999n 0.0 0.3333333333333333 0.6666666666666666 0.3333333333333333 0.4444444444444444
2190n 0.6666666666666666 0.0 0.3333333333333333 0.6666666666666666 0.7777777777777778
2199.999n 0.6666666666666666 0.0 0.3333333333333333 0.6666666666666666 0.7777777777777778
2200n 1.0 1.0 0.3333333333333333 1.0 1.7777777777777777
2209.999n 1.0 1.0 0.3333333333333333 1.0 1.7777777777777777
2210n 0.0 1.0 1.0 1.0 1.0
2219.999n 0.0 1.0 1.0 1.0 1.0
2220n 0.0 0.6666666666666666 1.0 0.3333333333333333 0.7777777777777778
2229.999n 0.0 0.6666666666666666 1.0 0.3333333333333333 0.7777777777777778
2230n 0.6666666666666666 1.0 0.0 1.0 1.3333333333333333
2239.999n 0.6666666666666666 1.0 0.0 1.0 1.3333333333333333
2240n 0.6666666666666666 0.6666666666666666 1.0 1.0 1.4444444444444444
2249.999n 0.6666666666666666 0.6666666666666666 1.0 1.0 1.4444444444444444
2250n 1.0 1.0 0.0 1.0 1.6666666666666667
2259.999n 1.0 1.0 0.0 1.0 1.6666666666666667
2260n 0.0 0.6666666666666666 0.0 0.0 0.4444444444444444
2269.999n 0.0 0.6666666666666666 0.0 0.0 0.4444444444444444
2270n 1.0 0.3333333333333333 0.6666666666666666 1.0 1.4444444444444444
2279.999n 1.0 0.3333333333333333 0.6666666666666666 1.0 1.4444444444444444
2280n 1.0 0.6666666666666666 0.6666666666666666 0.0 1.6666666666666667
2289.999n 1.0 0.6666666666666666 0.6666666666666666 0.0 1.6666666666666667
2290n 1.0 0.0 1.0 0.3333333333333333 1.3333333333333333
2299.999n 1.0 0.0 1.0 0.3333333333333333 1.3333333333333333
2300n 0.0 0.0 0.6666666666666666 1.0 0.2222222222222222
2309.999n 0.0 0.0 0.6666666666666666 1.0 0.2222222222222222
2310n 0.6666666666666666 0.3333333333333333 0.0 0.6666666666666666 0.8888888888888888
2319.999n 0.6666666666666666 0.3333333333333333 0.0 0.6666666666666666 0.8888888888888888
2320n 0.6666666666666666 1.0 0.6666666666666666 0.6666666666666666 1.5555555555555556
2329.999n 0.6666666666666666 1.0 0.6666666666666666 0.6666666666666666 1.5555555555555556
2330n 1.0 0.0 0.6666666666666666 1.0 1.2222222222222223
2339.999n 1.0 0.0 0.6666666666666666 1.0 1.2222222222222223
2340n 1.0 0.0 1.0 0.3333333333333333 1.3333333333333333
2349.999n 1.0 0.0 1.0 0.3333333333333333 1.3333333333333333
2350n 1.0 1.0 0.3333333333333333 0.3333333333333333 1.7777777777777777
2359.999n 1.0 1.0 0.3333333333333333 0.3333333333333333 1.7777777777777777
2360n 0.3333333333333333 1.0 0.0 1.0 1.0
2369.999n 0.3333333333333333 1.0 0.0 1.0 1.0
2370n 0.6666666666666666 0.3333333333333333 0.3333333333333333 1.0 1.0
2379.999n 0.6666666666666666 0.3333333333333333 0.3333333333333333 1.0 1.0
2380n 0.3333333333333333 0.0 0.3333333333333333 0.3333333333333333 0.4444444444444444
2389.999n 0.3333333333333333 0.0 0.3333333333333333 0.3333333333333333 0.4444444444444444
2390n 0.3333333333333333 0.3333333333333333 0.0 0.0 0.5555555555555556
2399.999n 0.3333333333333333 0.3333333333333333 0.0 0.0 0.5555555555555556
2400n 0.6666666666666666 0.3333333333333333 0.3333333333333333 0.6666666666666666 1.0
2409.999n 0.6666666666666666 0.3333333333333333 0.3333333333333333 0.6666666666666666 1.0
2410n 0.0 0.0 0.6666666666666666 0.0 0.2222222222222222
2419.999n 0.0 0.0 0.6666666666666666 0.0 0.2222222222222222
2420n 0.0 0.3333333333333333 0.3333333333333333 0.3333333333333333 0.3333333333333333
2429.999n 0.0 0.3333333333333333 0.3333333333333333 0.3333333333333333 0.3333333333333333
2430n 0.3333333333333333 0.6666666666666666 0.0 0.3333333333333333 0.7777777777777778
2439.999n 0.3333333333333333 0.6666666666666666 0.0 0.3333333333333333 0.7777777777777778
2440n 0.0 0.6666666666666666 1.0 0.0 0.7777777777777778
2449.999n 0.0 0.6666666666666666 1.0 0.0 0.7777777777777778
2450n 1.0 1.0 0.6666666666666666 0.0 1.8888888888888888
2459.999n 1.0 1.0 0.6666666666666666 0.0 1.8888888888888888
2460n 0.3333333333333333 1.0 1.0 0.0 1.3333333333333333
2469.999n 0.3333333333333333 1.0 1.0 0.0 1.3333333333333333
2470n 0.6666666666666666 0.6666666666666666 0.6666666666666666 1.0 1.3333333333333333
2479.999n 0.6666666666666666 0.6666666666666666 0.6666666666666666 1.0 1.3333333333333333
2480n 0.3333333333333333 1.0 0.0 0.6666666666666666 1.0
2489.999n 0.3333333333333333 1.0 0.0 0.6666666666666666 1.0
2490n 0.6666666666666666 1.0 0.0 0.3333333333333333 1.3333333333333333
2499.999n 0.6666666666666666 1.0 0.0 0.3333333333333333 1.3333333333333333
2500n 1.0 0.0 0.0 0.3333333333333333 1.0
2509.999n 1.0 0.0 0.0 0.3333333333333333 1.0
2510n 0.6666666666666666 1.0 0.3333333333333333 0.0 1.4444444444444444
2519.999n 0.6666666666666666 1.0 0.3333333333333333 0.0 1.4444444444444444
2520n 0.6666666666666666 0.6666666666666666 0.6666666666666666 1.0 1.3333333333333333
2529.999n 0.6666666666666666 0.6666666666666666 0.6666666666666666 1.0 1.3333333333333333
2530n 0.0 0.3333333333333333 0.6666666666666666 0.0 0.4444444444444444
2539.999n 0.0 0.3333333333333333 0.6666666666666666 0.0 0.4444444444444444
2540n 0.3333333333333333 0.6666666666666666 1.0 0.6666666666666666 1.1111111111111112
2549.999n 0.3333333333333333 0.6666666666666666 1.0 0.6666666666666666 1.1111111111111112
2550n 1.0 0.0 0.6666666666666666 0.3333333333333333 1.2222222222222223
2559.999n 1.0 0.0 0.6666666666666666 0.3333333333333333 1.2222222222222223
2560n 0.6666666666666666 0.0 1.0 0.3333333333333333 1.0
2569.999n 0.6666666666666666 0.0 1.0 0.3333333333333333 1.0
2570n 0.3333333333333333 0.3333333333333333 0.3333333333333333 0.3333333333333333 0.6666666666666666
2579.999n 0.3333333333333333 0.3333333333333333 0.3333333333333333 0.3333333333333333 0.6666666666666666
2580n 1.0 0.6666666666666666 1.0 0.6666666666666666 1.7777777777777777
2589.999n 1.0 0.6666666666666666 1.0 0.6666666666666666 1.7777777777777777
2590n 0.3333333333333333 0.0 0.3333333333333333 0.3333333333333333 0.4444444444444444
2599.999n 0.3333333333333333 0.0 0.3333333333333333 0.3333333333333333 0.4444444444444444
2600n 0.0 0.6666666666666666 1.0 0.6666666666666666 0.7777777777777778
2609.999n 0.0 0.6666666666666666 1.0 0.6666666666666666 0.7777777777777778
2610n 0.0 1.0 0.6666666666666666 0.6666666666666666 0.8888888888888888
2619.999n 0.0 1.0 0.6666666666666666 0.6666666666666666 0.8888888888888888
2620n 0.6666666666666666 0.6666666666666666 0.3333333333333333 0.0 1.2222222222222223
2629.999n 0.6666666666666666 0.6666666666666666 0.3333333333333333 0.0 1.2222222222222223
2630n 0.6666666666666666 0.0 1.0 0.3333333333333333 1.0
2639.999n 0.6666666666666666 0.0 1.0 0.3333333333333333 1.0
2640n 0.0 0.3333333333333333 0.6666666666666666 0.6666666666666666 0.4444444444444444
2649.999n 0.0 0.3333333333333333 0.6666666666666666 0.6666666666666666 0.4444444444444444
2650n 1.0 0.3333333333333333 1.0 0.0 1.5555555555555556
2659.999n 1.0 0.3333333333333333 1.0 0.0 1.5555555555555556
2660n 1.0 0.6666666666666666 0.0 0.0 1.4444444444444444
2669.999n 1.0 0.6666666666666666 0.0 0.0 1.4444444444444444
2670n 1.0 0.3333333333333333 0.3333333333333333 0.3333333333333333 1.3333333333333333
2679.999n 1.0 0.3333333333333333 0.3333333333333333 0.3333333333333333 1.3333333333333333
2680n 0.6666666666666666 0.0 1.0 1.0 1.0
2689.999n 0.6666666666666666 0.0 1.0 1.0 1.0
2690n 0.0 1.0 0.3333333333333333 0.0 0.7777777777777778
2699.999n 0.0 1.0 0.3333333333333333 0.0 0.7777777777777778
2700n 0.0 0.3333333333333333 0.6666666666666666 0.3333333333333333 0.4444444444444444
2709.999n 0.0 0.3333333333333333 0.6666666666666666 0.3333333333333333 0.4444444444444444
2710n 0.6666666666666666 0.6666666666666666 0.3333333333333333 0.6666666666666666 1.2222222222222223
2719.999n 0.6666666666666666 0.6666666666666666 0.3333333333333333 0.6666666666666666 1.2222222222222223
2720n 0.0 0.3333333333333333 0.0 0.6666666666666666 0.2222222222222222
2729.999n 0.0 0.3333333333333333 0.0 0.6666666666666666 0.2222222222222222
2730n 0.0 0.3333333333333333 1.0 0.6666666666666666 0.5555555555555556
2739.999n 0.0 0.3333333333333333 1.0 0.6666666666666666 0.5555555555555556
2740n 0.0 0.6666666666666666 0.6666666666666666 1.0 0.6666666666666666
2749.999n 0.0 0.6666666666666666 0.6666666666666666 1.0 0.6666666666666666
2750n 0.6666666666666666 1.0 1.0 0.6666666666666666 1.6666666666666667
2759.999n 0.6666666666666666 1.0 1.0 0.6666666666666666 1.6666666666666667
2760n 0.0 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.5555555555555556
2769.999n 0.0 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.5555555555555556
2770n 0.3333333333333333 0.3333333333333333 0.0 0.6666666666666666 0.5555555555555556
2779.999n 0.3333333333333333 0.3333333333333333 0.0 0.6666666666666666 0.5555555555555556
2780n 0.3333333333333333 1.0 1.0 0.0 1.3333333333333333
2789.999n 0.3333333333333333 1.0 1.0 0.0 1.3333333333333333
2790n 0.3333333333333333 0.3333333333333333 0.6666666666666666 0.6666666666666666 0.7777777777777778
2799.999n 0.3333333333333333 0.3333333333333333 0.6666666666666666 0.6666666666666666 0.7777777777777778
2800n 0.6666666666666666 1.0 0.0 0.0 1.3333333333333333
2809.999n 0.6666666666666666 1.0 0.0 0.0 1.3333333333333333
2810n 0.0 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.5555555555555556
2819.999n 0.0 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.5555555555555556
2820n 0.3333333333333333 0.6666666666666666 1.0 0.0 1.1111111111111112
2829.999n 0.3333333333333333 0.6666666666666666 1.0 0.0 1.1111111111111112
2830n 1.0 1.0 0.3333333333333333 0.0 1.7777777777777777
2839.999n 1.0 1.0 0.3333333333333333 0.0 1.7777777777777777
2840n 0.6666666666666666 0.6666666666666666 1.0 0.0 1.4444444444444444
2849.999n 0.6666666666666666 0.6666666666666666 1.0 0.0 1.4444444444444444
2850n 0.6666666666666666 0.3333333333333333 0.3333333333333333 0.6666666666666666 1.0
2859.999n 0.6666666666666666 0.3333333333333333 0.3333333333333333 0.6666666666666666 1.0
2860n 0.3333333333333333 1.0 0.0 0.0 1.0
2869.999n 0.3333333333333333 1.0 0.0 0.0 1.0
2870n 1.0 0.3333333333333333 0.6666666666666666 0.0 1.4444444444444444
2879.999n 1.0 0.3333333333333333 0.6666666666666666 0.0 1.4444444444444444
2880n 1.0 0.6666666666666666 1.0 1.0 1.7777777777777777
2889.999n 1.0 0.6666666666666666 1.0 1.0 1.7777777777777777
2890n 0.3333333333333333 0.3333333333333333 0.0 0.0 0.5555555555555556
2899.999n 0.3333333333333333 0.3333333333333333 0.0 0.0 0.5555555555555556
2900n 0.3333333333333333 1.0 1.0 0.3333333333333333 1.3333333333333333
2909.999n 0.3333333333333333 1.0 1.0 0.3333333333333333 1.3333333333333333
2910n 0.3333333333333333 1.0 0.3333333333333333 0.6666666666666666 1.1111111111111112
2919.999n 0.3333333333333333 1.0 0.3333333333333333 0.6666666666666666 1.1111111111111112
2920n 0.3333333333333333 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.8888888888888888
2929.999n 0.3333333333333333 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.8888888888888888
2930n 1.0 0.3333333333333333 0.6666666666666666 1.0 1.4444444444444444
2939.999n 1.0 0.3333333333333333 0.6666666666666666 1.0 1.4444444444444444
2940n 1.0 1.0 0.6666666666666666 1.0 1.8888888888888888
2949.999n 1.0 1.0 0.6666666666666666 1.0 1.8888888888888888
2950n 1.0 0.0 0.6666666666666666 0.3333333333333333 1.2222222222222223
2959.999n 1.0 0.0 0.6666666666666666 0.3333333333333333 1.2222222222222223
2960n 1.0 0.3333333333333333 1.0 0.0 1.5555555555555556
2969.999n 1.0 0.3333333333333333 1.0 0.0 1.5555555555555556
2970n 0.3333333333333333 1.0 0.3333333333333333 1.0 1.1111111111111112
2979.999n 0.3333333333333333 1.0 0.3333333333333333 1.0 1.1111111111111112
2980n 0.6666666666666666 0.3333333333333333 0.3333333333333333 0.0 1.0
2989.999n 0.6666666666666666 0.3333333333333333 0.3333333333333333 0.0 1.0
2990n 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.6666666666666666 1.1111111111111112
2999.999n 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.6666666666666666 1.1111111111111112
3000n 0.0 0.0 1.0 0.6666666666666666 0.3333333333333333
3009.999n 0.0 0.0 1.0 0.6666666666666666 0.3333333333333333
3010n 0.3333333333333333 0.3333333333333333 0.0 0.6666666666666666 0.5555555555555556
3019.999n 0.3333333333333333 0.3333333333333333 0.0 0.6666666666666666 0.5555555555555556
3020n 0.6666666666666666 1.0 0.6666666666666666 1.0 1.5555555555555556
3029.999n 0.6666666666666666 1.0 0.6666666666666666 1.0 1.5555555555555556
3030n 0.3333333333333333 0.0 0.0 0.3333333333333333 0.3333333333333333
3039.999n 0.3333333333333333 0.0 0.0 0.3333333333333333 0.3333333333333333
3040n 0.6666666666666666 1.0 0.3333333333333333 0.6666666666666666 1.4444444444444444
3049.999n 0.6666666666666666 1.0 0.3333333333333333 0.6666666666666666 1.4444444444444444
3050n 1.0 0.6666666666666666 0.0 1.0 1.4444444444444444
3059.999n 1.0 0.6666666666666666 0.0 1.0 1.4444444444444444
3060n 0.0 1.0 0.6666666666666666 0.3333333333333333 0.8888888888888888
3069.999n 0.0 1.0 0.6666666666666666 0.3333333333333333 0.8888888888888888
3070n 0.3333333333333333 1.0 0.0 0.3333333333333333 1.0
3079.999n 0.3333333333333333 1.0 0.0 0.3333333333333333 1.0
3080n 0.6666666666666666 0.6666666666666666 0.0 0.3333333333333333 1.1111111111111112
3089.999n 0.6666666666666666 0.6666666666666666 0.0 0.3333333333333333 1.1111111111111112
3090n 0.6666666666666666 1.0 1.0 1.0 1.6666666666666667
3099.999n 0.6666666666666666 1.0 1.0 1.0 1.6666666666666667
3100n 1.0 0.3333333333333333 0.3333333333333333 0.0 1.3333333333333333
3109.999n 1.0 0.3333333333333333 0.3333333333333333 0.0 1.3333333333333333
3110n 0.3333333333333333 0.0 0.0 0.6666666666666666 0.3333333333333333
3119.999n 0.3333333333333333 0.0 0.0 0.6666666666666666 0.3333333333333333
3120n 0.3333333333333333 0.6666666666666666 0.3333333333333333 1.0 0.8888888888888888
3129.999n 0.3333333333333333 0.6666666666666666 0.3333333333333333 1.0 0.8888888888888888
3130n 1.0 1.0 0.0 1.0 1.6666666666666667
3139.999n 1.0 1.0 0.0 1.0 1.6666666666666667
3140n 1.0 0.6666666666666666 0.3333333333333333 0.3333333333333333 1.5555555555555556
3149.999n 1.0 0.6666666666666666 0.3333333333333333 0.3333333333333333 1.5555555555555556
3150n 0.0 1.0 0.0 0.0 0.6666666666666666
3159.999n 0.0 1.0 0.0 0.0 0.6666666666666666
3160n 0.0 0.0 0.6666666666666666 0.6666666666666666 0.2222222222222222
3169.999n 0.0 0.0 0.6666666666666666 0.6666666666666666 0.2222222222222222
3170n 1.0 1.0 0.3333333333333333 1.0 1.7777777777777777
3179.999n 1.0 1.0 0.3333333333333333 1.0 1.7777777777777777
3180n 1.0 0.3333333333333333 0.6666666666666666 0.0 1.4444444444444444
3189.999n 1.0 0.3333333333333333 0.6666666666666666 0.0 1.4444444444444444
3190n 0.0 0.3333333333333333 1.0 1.0 0.5555555555555556
3199.999n 0.0 0.3333333333333333 1.0 1.0 0.5555555555555556
3200n 0.6666666666666666 0.3333333333333333 0.3333333333333333 1.0 1.0
3209.999n 0.6666666666666666 0.3333333333333333 0.3333333333333333 1.0 1.0
3210n 0.0 1.0 0.3333333333333333 0.3333333333333333 0.7777777777777778
3219.999n 0.0 1.0 0.3333333333333333 0.3333333333333333 0.7777777777777778
3220n 0.6666666666666666 0.0 1.0 0.0 1.0
3229.999n 0.6666666666666666 0.0 1.0 0.0 1.0
3230n 1.0 0.3333333333333333 0.0 1.0 1.2222222222222223
3239.999n 1.0 0.3333333333333333 0.0 1.0 1.2222222222222223
3240n 1.0 0.3333333333333333 0.0 0.6666666666666666 1.2222222222222223
3249.999n 1.0 0.3333333333333333 0.0 0.6666666666666666 1.2222222222222223
3250n 0.3333333333333333 0.6666666666666666 1.0 0.0 1.1111111111111112
3259.999n 0.3333333333333333 0.6666666666666666 1.0 0.0 1.1111111111111112
3260n 0.3333333333333333 0.0 0.3333333333333333 0.6666666666666666 0.4444444444444444
3269.999n 0.3333333333333333 0.0 0.3333333333333333 0.6666666666666666 0.4444444444444444
3270n 0.3333333333333333 1.0 1.0 0.3333333333333333 1.3333333333333333
3279.999n 0.3333333333333333 1.0 1.0 0.3333333333333333 1.3333333333333333
3280n 0.0 1.0 0.6666666666666666 0.3333333333333333 0.8888888888888888
3289.999n 0.0 1.0 0.6666666666666666 0.3333333333333333 0.8888888888888888
3290n 1.0 1.0 0.6666666666666666 0.3333333333333333 1.8888888888888888
3299.999n 1.0 1.0 0.6666666666666666 0.3333333333333333 1.8888888888888888
3300n 0.3333333333333333 0.3333333333333333 0.0 0.0 0.5555555555555556
3309.999n 0.3333333333333333 0.3333333333333333 0.0 0.0 0.5555555555555556
3310n 1.0 1.0 0.6666666666666666 0.6666666666666666 1.8888888888888888
3319.999n 1.0 1.0 0.6666666666666666 0.6666666666666666 1.8888888888888888
3320n 0.6666666666666666 0.0 0.6666666666666666 1.0 0.8888888888888888
3329.999n 0.6666666666666666 0.0 0.6666666666666666 1.0 0.8888888888888888
3330n 0.6666666666666666 0.6666666666666666 0.3333333333333333 0.3333333333333333 1.2222222222222223
3339.999n 0.6666666666666666 0.6666666666666666 0.3333333333333333 0.3333333333333333 1.2222222222222223
3340n 0.6666666666666666 0.6666666666666666 0.6666666666666666 1.0 1.3333333333333333
3349.999n 0.6666666666666666 0.6666666666666666 0.6666666666666666 1.0 1.3333333333333333
3350n 0.0 0.3333333333333333 1.0 0.3333333333333333 0.5555555555555556
3359.999n 0.0 0.3333333333333333 1.0 0.3333333333333333 0.5555555555555556
3360n 1.0 1.0 0.3333333333333333 0.6666666666666666 1.7777777777777777
3369.999n 1.0 1.0 0.3333333333333333 0.6666666666666666 1.7777777777777777
3370n 1.0 0.3333333333333333 0.0 0.6666666666666666 1.2222222222222223
3379.999n 1.0 0.3333333333333333 0.0 0.6666666666666666 1.2222222222222223
3380n 0.0 0.0 0.3333333333333333 0.3333333333333333 0.1111111111111111
3389.999n 0.0 0.0 0.3333333333333333 0.3333333333333333 0.1111111111111111
3390n 0.0 0.0 0.3333333333333333 1.0 0.1111111111111111
3399.999n 0.0 0.0 0.3333333333333333 1.0 0.1111111111111111
3400n 0.6666666666666666 0.6666666666666666 0.3333333333333333 1.0 1.2222222222222223
3409.999n 0.6666666666666666 0.6666666666666666 0.3333333333333333 1.0 1.2222222222222223
3410n 0.0 1.0 0.3333333333333333 1.0 0.7777777777777778
3419.999n 0.0 1.0 0.3333333333333333 1.0 0.7777777777777778
3420n 1.0 0.3333333333333333 0.3333333333333333 1.0 1.3333333333333333
3429.999n 1.0 0.3333333333333333 0.3333333333333333 1.0 1.3333333333333333
3430n 1.0 0.3333333333333333 0.0 0.0 1.2222222222222223
3439.999n 1.0 0.3333333333333333 0.0 0.0 1.2222222222222223
3440n 0.6666666666666666 0.0 1.0 0.6666666666666666 1.0
3449.999n 0.6666666666666666 0.0 1.0 0.6666666666666666 1.0
3450n 0.0 0.6666666666666666 0.3333333333333333 1.0 0.5555555555555556
3459.999n 0.0 0.6666666666666666 0.3333333333333333 1.0 0.5555555555555556
3460n 0.3333333333333333 0.6666666666666666 1.0 1.0 1.1111111111111112
3469.999n 0.3333333333333333 0.6666666666666666 1.0 1.0 1.1111111111111112
3470n 0.6666666666666666 0.0 0.6666666666666666 0.6666666666666666 0.8888888888888888
3479.999n 0.6666666666666666 0.0 0.6666666666666666 0.6666666666666666 0.8888888888888888
3480n 0.3333333333333333 0.6666666666666666 1.0 0.6666666666666666 1.1111111111111112
3489.999n 0.3333333333333333 0.6666666666666666 1.0 0.6666666666666666 1.1111111111111112
3490n 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.3333333333333333 1.1111111111111112
3499.999n 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.3333333333333333 1.1111111111111112
3500n 1.0 1.0 0.6666666666666666 0.0 1.8888888888888888
3509.999n 1.0 1.0 0.6666666666666666 0.0 1.8888888888888888
3510n 0.6666666666666666 0.3333333333333333 0.3333333333333333 0.0 1.0
3519.999n 0.6666666666666666 0.3333333333333333 0.3333333333333333 0.0 1.0
3520n 0.3333333333333333 0.3333333333333333 0.6666666666666666 1.0 0.7777777777777778
3529.999n 0.3333333333333333 0.3333333333333333 0.6666666666666666 1.0 0.7777777777777778
3530n 1.0 0.0 0.3333333333333333 1.0 1.1111111111111112
3539.999n 1.0 0.0 0.3333333333333333 1.0 1.1111111111111112
3540n 1.0 0.3333333333333333 0.6666666666666666 1.0 1.4444444444444444
3549.999n 1.0 0.3333333333333333 0.6666666666666666 1.0 1.4444444444444444
3550n 0.3333333333333333 1.0 0.0 0.0 1.0
3559.999n 0.3333333333333333 1.0 0.0 0.0 1.0
3560n 0.6666666666666666 1.0 0.6666666666666666 0.0 1.5555555555555556
3569.999n 0.6666666666666666 1.0 0.6666666666666666 0.0 1.5555555555555556
3570n 0.6666666666666666 1.0 1.0 1.0 1.6666666666666667
3579.999n 0.6666666666666666 1.0 1.0 1.0 1.6666666666666667
3580n 0.6666666666666666 0.3333333333333333 0.3333333333333333 0.0 1.0
3589.999n 0.6666666666666666 0.3333333333333333 0.3333333333333333 0.0 1.0
3590n 0.0 0.6666666666666666 0.0 0.3333333333333333 0.4444444444444444
3599.999n 0.0 0.6666666666666666 0.0 0.3333333333333333 0.4444444444444444
3600n 1.0 0.3333333333333333 0.6666666666666666 1.0 1.4444444444444444
3609.999n 1.0 0.3333333333333333 0.6666666666666666 1.0 1.4444444444444444
3610n 1.0 0.6666666666666666 0.6666666666666666 0.3333333333333333 1.6666666666666667
3619.999n 1.0 0.6666666666666666 0.6666666666666666 0.3333333333333333 1.6666666666666667
3620n 1.0 0.0 0.3333333333333333 0.0 1.1111111111111112
3629.999n 1.0 0.0 0.3333333333333333 0.0 1.1111111111111112
3630n 1.0 0.0 0.6666666666666666 0.0 1.2222222222222223
3639.999n 1.0 0.0 0.6666666666666666 0.0 1.2222222222222223
3640n 0.3333333333333333 1.0 0.3333333333333333 0.3333333333333333 1.1111111111111112
3649.999n 0.3333333333333333 1.0 0.3333333333333333 0.3333333333333333 1.1111111111111112
3650n 0.6666666666666666 0.3333333333333333 1.0 1.0 1.2222222222222223
3659.999n 0.6666666666666666 0.3333333333333333 1.0 1.0 1.2222222222222223
3660n 0.0 0.0 0.0 0.6666666666666666 0.0
3669.999n 0.0 0.0 0.0 0.6666666666666666 0.0
3670n 0.6666666666666666 0.0 0.3333333333333333 0.3333333333333333 0.7777777777777778
3679.999n 0.6666666666666666 0.0 0.3333333333333333 0.3333333333333333 0.7777777777777778
3680n 0.6666666666666666 0.3333333333333333 0.0 0.6666666666666666 0.8888888888888888
3689.999n 0.6666666666666666 0.3333333333333333 0.0 0.6666666666666666 0.8888888888888888
3690n 0.6666666666666666 1.0 0.3333333333333333 0.6666666666666666 1.4444444444444444
3699.999n 0.6666666666666666 1.0 0.3333333333333333 0.6666666666666666 1.4444444444444444
3700n 0.6666666666666666 0.6666666666666666 0.3333333333333333 0.0 1.2222222222222223
3709.999n 0.6666666666666666 0.6666666666666666 0.3333333333333333 0.0 1.2222222222222223
3710n 1.0 1.0 0.3333333333333333 0.6666666666666666 1.7777777777777777
3719.999n 1.0 1.0 0.3333333333333333 0.6666666666666666 1.7777777777777777
3720n 0.3333333333333333 0.6666666666666666 1.0 0.0 1.1111111111111112
3729.999n 0.3333333333333333 0.6666666666666666 1.0 0.0 1.1111111111111112
3730n 0.0 0.6666666666666666 0.3333333333333333 0.3333333333333333 0.5555555555555556
3739.999n 0.0 0.6666666666666666 0.3333333333333333 0.3333333333333333 0.5555555555555556
3740n 1.0 0.0 0.6666666666666666 1.0 1.2222222222222223
3749.999n 1.0 0.0 0.6666666666666666 1.0 1.2222222222222223
3750n 0.3333333333333333 0.3333333333333333 1.0 1.0 0.8888888888888888
3759.999n 0.3333333333333333 0.3333333333333333 1.0 1.0 0.8888888888888888
3760n 1.0 0.3333333333333333 0.6666666666666666 0.6666666666666666 1.4444444444444444
3769.999n 1.0 0.3333333333333333 0.6666666666666666 0.6666666666666666 1.4444444444444444
3770n 0.3333333333333333 1.0 0.0 0.0 1.0
3779.999n 0.3333333333333333 1.0 0.0 0.0 1.0
3780n 0.6666666666666666 0.3333333333333333 0.6666666666666666 1.0 1.1111111111111112
3789.999n 0.6666666666666666 0.3333333333333333 0.6666666666666666 1.0 1.1111111111111112
3790n 0.0 0.6666666666666666 0.0 0.3333333333333333 0.4444444444444444
3799.999n 0.0 0.6666666666666666 0.0 0.3333333333333333 0.4444444444444444
3800n 1.0 0.6666666666666666 1.0 0.6666666666666666 1.7777777777777777
3809.999n 1.0 0.6666666666666666 1.0 0.6666666666666666 1.7777777777777777
3810n 0.0 0.3333333333333333 0.3333333333333333 0.3333333333333333 0.3333333333333333
3819.999n 0.0 0.3333333333333333 0.3333333333333333 0.3333333333333333 0.3333333333333333
3820n 1.0 1.0 0.0 0.3333333333333333 1.6666666666666667
3829.999n 1.0 1.0 0.0 0.3333333333333333 1.6666666666666667
3830n 1.0 0.0 1.0 1.0 1.3333333333333333
3839.999n 1.0 0.0 1.0 1.0 1.3333333333333333
3840n 0.3333333333333333 1.0 1.0 0.3333333333333333 1.3333333333333333
3849.999n 0.3333333333333333 1.0 1.0 0.3333333333333333 1.3333333333333333
3850n 0.6666666666666666 0.6666666666666666 0.6666666666666666 0.3333333333333333 1.3333333333333333
3859.999n 0.6666666666666666 0.6666666666666666 0.6666666666666666 0.3333333333333333 1.3333333333333333
3860n 0.3333333333333333 0.6666666666666666 0.0 0.0 0.7777777777777778
3869.999n 0.3333333333333333 0.6666666666666666 0.0 0.0 0.7777777777777778
3870n 0.3333333333333333 1.0 0.0 0.3333333333333333 1.0
3879.999n 0.3333333333333333 1.0 0.0 0.3333333333333333 1.0
3880n 1.0 1.0 0.6666666666666666 1.0 1.8888888888888888
3889.999n 1.0 1.0 0.6666666666666666 1.0 1.8888888888888888
3890n 1.0 0.3333333333333333 0.3333333333333333 0.6666666666666666 1.3333333333333333
3899.999n 1.0 0.3333333333333333 0.3333333333333333 0.6666666666666666 1.3333333333333333
3900n 0.6666666666666666 0.0 0.3333333333333333 1.0 0.7777777777777778
3909.999n 0.6666666666666666 0.0 0.3333333333333333 1.0 0.7777777777777778
3910n 0.3333333333333333 0.0 0.6666666666666666 0.3333333333333333 0.5555555555555556
3919.999n 0.3333333333333333 0.0 0.6666666666666666 0.3333333333333333 0.5555555555555556
3920n 0.0 0.0 0.6666666666666666 0.3333333333333333 0.2222222222222222
3929.999n 0.0 0.0 0.6666666666666666 0.3333333333333333 0.2222222222222222
3930n 1.0 0.0 1.0 0.3333333333333333 1.3333333333333333
3939.999n 1.0 0.0 1.0 0.3333333333333333 1.3333333333333333
3940n 0.0 1.0 0.3333333333333333 0.3333333333333333 0.7777777777777778
3949.999n 0.0 1.0 0.3333333333333333 0.3333333333333333 0.7777777777777778
3950n 0.0 1.0 0.3333333333333333 0.3333333333333333 0.7777777777777778
3959.999n 0.0 1.0 0.3333333333333333 0.3333333333333333 0.7777777777777778
3960n 0.0 0.6666666666666666 0.6666666666666666 0.0 0.6666666666666666
3969.999n 0.0 0.6666666666666666 0.6666666666666666 0.0 0.6666666666666666
3970n 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.6666666666666666 1.1111111111111112
3979.999n 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.6666666666666666 1.1111111111111112
3980n 0.3333333333333333 1.0 0.6666666666666666 0.0 1.2222222222222223
3989.999n 0.3333333333333333 1.0 0.6666666666666666 0.0 1.2222222222222223
3990n 0.0 1.0 0.6666666666666666 0.3333333333333333 0.8888888888888888
3999.999n 0.0 1.0 0.6666666666666666 0.3333333333333333 0.8888888888888888
4000n 1.0 0.6666666666666666 0.6666666666666666 1.0 1.6666666666666667
4009.999n 1.0 0.6666666666666666 0.6666666666666666 1.0 1.6666666666666667
4010n 0.3333333333333333 0.6666666666666666 0.3333333333333333 0.0 0.8888888888888888
4019.999n 0.3333333333333333 0.6666666666666666 0.3333333333333333 0.0 0.8888888888888888
4020n 0.6666666666666666 0.6666666666666666 1.0 0.0 1.4444444444444444
4029.999n 0.6666666666666666 0.6666666666666666 1.0 0.0 1.4444444444444444
4030n 0.0 1.0 0.0 1.0 0.6666666666666666
4039.999n 0.0 1.0 0.0 1.0 0.6666666666666666
4040n 1.0 1.0 0.0 1.0 1.6666666666666667
4049.999n 1.0 1.0 0.0 1.0 1.6666666666666667
4050n 0.6666666666666666 0.6666666666666666 0.3333333333333333 0.3333333333333333 1.2222222222222223
4059.999n 0.6666666666666666 0.6666666666666666 0.3333333333333333 0.3333333333333333 1.2222222222222223
4060n 1.0 1.0 0.0 0.0 1.6666666666666667
4069.999n 1.0 1.0 0.0 0.0 1.6666666666666667
4070n 0.6666666666666666 0.6666666666666666 0.6666666666666666 0.3333333333333333 1.3333333333333333
4079.999n 0.6666666666666666 0.6666666666666666 0.6666666666666666 0.3333333333333333 1.3333333333333333
4080n 0.0 0.0 0.6666666666666666 0.6666666666666666 0.2222222222222222
4089.999n 0.0 0.0 0.6666666666666666 0.6666666666666666 0.2222222222222222
4090n 0.6666666666666666 0.6666666666666666 1.0 0.6666666666666666 1.4444444444444444
4099.999n 0.6666666666666666 0.6666666666666666 1.0 0.6666666666666666 1.4444444444444444
4100n 0.6666666666666666 1.0 0.0 0.6666666666666666 1.3333333333333333
4109.999n 0.6666666666666666 1.0 0.0 0.6666666666666666 1.3333333333333333
4110n 0.0 0.0 0.3333333333333333 0.3333333333333333 0.1111111111111111
4119.999n 0.0 0.0 0.3333333333333333 0.3333333333333333 0.1111111111111111
4120n 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.0 1.1111111111111112
4129.999n 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.0 1.1111111111111112
4130n 0.0 0.3333333333333333 0.3333333333333333 0.6666666666666666 0.3333333333333333
4139.999n 0.0 0.3333333333333333 0.3333333333333333 0.6666666666666666 0.3333333333333333
4140n 0.0 0.6666666666666666 1.0 0.6666666666666666 0.7777777777777778
4149.999n 0.0 0.6666666666666666 1.0 0.6666666666666666 0.7777777777777778
4150n 0.3333333333333333 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.8888888888888888
4159.999n 0.3333333333333333 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.8888888888888888
4160n 0.3333333333333333 0.3333333333333333 0.0 0.3333333333333333 0.5555555555555556
4169.999n 0.3333333333333333 0.3333333333333333 0.0 0.3333333333333333 0.5555555555555556
4170n 1.0 0.0 0.3333333333333333 0.0 1.1111111111111112
4179.999n 1.0 0.0 0.3333333333333333 0.0 1.1111111111111112
4180n 0.6666666666666666 0.0 0.3333333333333333 0.3333333333333333 0.7777777777777778
4189.999n 0.6666666666666666 0.0 0.3333333333333333 0.3333333333333333 0.7777777777777778
4190n 1.0 0.6666666666666666 0.6666666666666666 0.0 1.6666666666666667
4199.999n 1.0 0.6666666666666666 0.6666666666666666 0.0 1.6666666666666667
4200n 0.6666666666666666 0.3333333333333333 0.3333333333333333 0.6666666666666666 1.0
4209.999n 0.6666666666666666 0.3333333333333333 0.3333333333333333 0.6666666666666666 1.0
4210n 0.0 0.6666666666666666 0.6666666666666666 1.0 0.6666666666666666
4219.999n 0.0 0.6666666666666666 0.6666666666666666 1.0 0.6666666666666666
4220n 0.0 1.0 0.6666666666666666 0.3333333333333333 0.8888888888888888
4229.999n 0.0 1.0 0.6666666666666666 0.3333333333333333 0.8888888888888888
4230n 1.0 0.3333333333333333 0.0 1.0 1.2222222222222223
4239.999n 1.0 0.3333333333333333 0.0 1.0 1.2222222222222223
4240n 0.0 1.0 1.0 0.3333333333333333 1.0
4249.999n 0.0 1.0 1.0 0.3333333333333333 1.0
4250n 1.0 0.3333333333333333 0.3333333333333333 0.3333333333333333 1.3333333333333333
4259.999n 1.0 0.3333333333333333 0.3333333333333333 0.3333333333333333 1.3333333333333333
4260n 0.3333333333333333 0.6666666666666666 0.0 0.0 0.7777777777777778
4269.999n 0.3333333333333333 0.6666666666666666 0.0 0.0 0.7777777777777778
4270n 1.0 0.0 1.0 1.0 1.3333333333333333
4279.999n 1.0 0.0 1.0 1.0 1.3333333333333333
4280n 0.3333333333333333 1.0 0.6666666666666666 0.3333333333333333 1.2222222222222223
4289.999n 0.3333333333333333 1.0 0.6666666666666666 0.3333333333333333 1.2222222222222223
4290n 0.3333333333333333 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.8888888888888888
4299.999n 0.3333333333333333 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.8888888888888888
4300n 0.6666666666666666 0.6666666666666666 1.0 0.3333333333333333 1.4444444444444444
4309.999n 0.6666666666666666 0.6666666666666666 1.0 0.3333333333333333 1.4444444444444444
4310n 1.0 0.0 0.3333333333333333 0.0 1.1111111111111112
4319.999n 1.0 0.0 0.3333333333333333 0.0 1.1111111111111112
4320n 1.0 0.3333333333333333 0.3333333333333333 0.6666666666666666 1.3333333333333333
4329.999n 1.0 0.3333333333333333 0.3333333333333333 0.6666666666666666 1.3333333333333333
4330n 1.0 0.3333333333333333 0.0 0.6666666666666666 1.2222222222222223
4339.999n 1.0 0.3333333333333333 0.0 0.6666666666666666 1.2222222222222223
4340n 1.0 0.6666666666666666 1.0 0.3333333333333333 1.7777777777777777
4349.999n 1.0 0.6666666666666666 1.0 0.3333333333333333 1.7777777777777777
4350n 0.6666666666666666 0.0 0.0 0.3333333333333333 0.6666666666666666
4359.999n 0.6666666666666666 0.0 0.0 0.3333333333333333 0.6666666666666666
4360n 0.0 0.0 0.3333333333333333 1.0 0.1111111111111111
4369.999n 0.0 0.0 0.3333333333333333 1.0 0.1111111111111111
4370n 0.0 0.3333333333333333 0.3333333333333333 1.0 0.3333333333333333
4379.999n 0.0 0.3333333333333333 0.3333333333333333 1.0 0.3333333333333333
4380n 0.3333333333333333 0.3333333333333333 0.3333333333333333 1.0 0.6666666666666666
4389.999n 0.3333333333333333 0.3333333333333333 0.3333333333333333 1.0 0.6666666666666666
4390n 0.0 0.0 0.0 0.3333333333333333 0.0
4399.999n 0.0 0.0 0.0 0.3333333333333333 0.0
4400n 0.6666666666666666 0.0 0.0 0.0 0.6666666666666666
4409.999n 0.6666666666666666 0.0 0.0 0.0 0.6666666666666666
4410n 0.0 0.0 0.0 0.6666666666666666 0.0
4419.999n 0.0 0.0 0.0 0.6666666666666666 0.0
4420n 0.6666666666666666 0.0 0.0 1.0 0.6666666666666666
4429.999n 0.6666666666666666 0.0 0.0 1.0 0.6666666666666666
4430n 0.6666666666666666 0.6666666666666666 0.6666666666666666 0.3333333333333333 1.3333333333333333
4439.999n 0.6666666666666666 0.6666666666666666 0.6666666666666666 0.3333333333333333 1.3333333333333333
4440n 0.3333333333333333 1.0 0.0 1.0 1.0
4449.999n 0.3333333333333333 1.0 0.0 1.0 1.0
4450n 0.6666666666666666 1.0 0.6666666666666666 0.3333333333333333 1.5555555555555556
4459.999n 0.6666666666666666 1.0 0.6666666666666666 0.3333333333333333 1.5555555555555556
4460n 0.3333333333333333 0.3333333333333333 1.0 0.3333333333333333 0.8888888888888888
4469.999n 0.3333333333333333 0.3333333333333333 1.0 0.3333333333333333 0.8888888888888888
4470n 0.3333333333333333 0.6666666666666666 0.6666666666666666 1.0 1.0
4479.999n 0.3333333333333333 0.6666666666666666 0.6666666666666666 1.0 1.0
4480n 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.3333333333333333 1.1111111111111112
4489.999n 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.3333333333333333 1.1111111111111112
4490n 0.3333333333333333 1.0 0.0 0.3333333333333333 1.0
4499.999n 0.3333333333333333 1.0 0.0 0.3333333333333333 1.0
4500n 1.0 0.6666666666666666 0.6666666666666666 0.3333333333333333 1.6666666666666667
4509.999n 1.0 0.6666666666666666 0.6666666666666666 0.3333333333333333 1.6666666666666667
4510n 0.6666666666666666 0.3333333333333333 1.0 0.0 1.2222222222222223
4519.999n 0.6666666666666666 0.3333333333333333 1.0 0.0 1.2222222222222223
4520n 0.3333333333333333 1.0 1.0 0.0 1.3333333333333333
4529.999n 0.3333333333333333 1.0 1.0 0.0 1.3333333333333333
4530n 0.3333333333333333 0.6666666666666666 0.0 0.3333333333333333 0.7777777777777778
4539.999n 0.3333333333333333 0.6666666666666666 0.0 0.3333333333333333 0.7777777777777778
4540n 1.0 0.0 0.6666666666666666 0.0 1.2222222222222223
4549.999n 1.0 0.0 0.6666666666666666 0.0 1.2222222222222223
4550n 0.0 0.3333333333333333 0.3333333333333333 0.6666666666666666 0.3333333333333333
4559.999n 0.0 0.3333333333333333 0.3333333333333333 0.6666666666666666 0.3333333333333333
4560n 0.3333333333333333 1.0 1.0 0.0 1.3333333333333333
4569.999n 0.3333333333333333 1.0 1.0 0.0 1.3333333333333333
4570n 0.0 0.3333333333333333 0.3333333333333333 0.3333333333333333 0.3333333333333333
4579.999n 0.0 0.3333333333333333 0.3333333333333333 0.3333333333333333 0.3333333333333333
4580n 0.6666666666666666 1.0 1.0 0.6666666666666666 1.6666666666666667
4589.999n 0.6666666666666666 1.0 1.0 0.6666666666666666 1.6666666666666667
4590n 1.0 1.0 0.6666666666666666 1.0 1.8888888888888888
4599.999n 1.0 1.0 0.6666666666666666 1.0 1.8888888888888888
4600n 0.6666666666666666 0.3333333333333333 0.3333333333333333 0.3333333333333333 1.0
4609.999n 0.6666666666666666 0.3333333333333333 0.3333333333333333 0.3333333333333333 1.0
4610n 0.3333333333333333 0.3333333333333333 0.3333333333333333 1.0 0.6666666666666666
4619.999n 0.3333333333333333 0.3333333333333333 0.3333333333333333 1.0 0.6666666666666666
4620n 0.0 1.0 0.0 0.0 0.6666666666666666
4629.999n 0.0 1.0 0.0 0.0 0.6666666666666666
4630n 0.3333333333333333 0.3333333333333333 0.3333333333333333 0.3333333333333333 0.6666666666666666
4639.999n 0.3333333333333333 0.3333333333333333 0.3333333333333333 0.3333333333333333 0.6666666666666666
4640n 0.6666666666666666 1.0 1.0 0.6666666666666666 1.6666666666666667
4649.999n 0.6666666666666666 1.0 1.0 0.6666666666666666 1.6666666666666667
4650n 0.6666666666666666 0.6666666666666666 1.0 1.0 1.4444444444444444
4659.999n 0.6666666666666666 0.6666666666666666 1.0 1.0 1.4444444444444444
4660n 0.0 0.0 1.0 0.3333333333333333 0.3333333333333333
4669.999n 0.0 0.0 1.0 0.3333333333333333 0.3333333333333333
4670n 0.6666666666666666 1.0 0.3333333333333333 0.0 1.4444444444444444
4679.999n 0.6666666666666666 1.0 0.3333333333333333 0.0 1.4444444444444444
4680n 1.0 0.3333333333333333 0.3333333333333333 0.3333333333333333 1.3333333333333333
4689.999n 1.0 0.3333333333333333 0.3333333333333333 0.3333333333333333 1.3333333333333333
4690n 0.3333333333333333 0.6666666666666666 0.0 0.6666666666666666 0.7777777777777778
4699.999n 0.3333333333333333 0.6666666666666666 0.0 0.6666666666666666 0.7777777777777778
4700n 0.6666666666666666 1.0 0.0 1.0 1.3333333333333333
4709.999n 0.6666666666666666 1.0 0.0 1.0 1.3333333333333333
4710n 0.3333333333333333 0.3333333333333333 1.0 0.0 0.8888888888888888
4719.999n 0.3333333333333333 0.3333333333333333 1.0 0.0 0.8888888888888888
4720n 0.3333333333333333 0.0 0.0 0.6666666666666666 0.3333333333333333
4729.999n 0.3333333333333333 0.0 0.0 0.6666666666666666 0.3333333333333333
4730n 0.0 0.3333333333333333 0.0 1.0 0.2222222222222222
4739.999n 0.0 0.3333333333333333 0.0 1.0 0.2222222222222222
4740n 1.0 0.6666666666666666 0.3333333333333333 0.0 1.5555555555555556
4749.999n 1.0 0.6666666666666666 0.3333333333333333 0.0 1.5555555555555556
4750n 1.0 0.6666666666666666 0.3333333333333333 1.0 1.5555555555555556
4759.999n 1.0 0.6666666666666666 0.3333333333333333 1.0 1.5555555555555556
4760n 0.3333333333333333 0.6666666666666666 1.0 0.0 1.1111111111111112
4769.999n 0.3333333333333333 0.6666666666666666 1.0 0.0 1.1111111111111112
4770n 1.0 1.0 0.3333333333333333 1.0 1.7777777777777777
4779.999n 1.0 1.0 0.3333333333333333 1.0 1.7777777777777777
4780n 1.0 0.0 1.0 0.3333333333333333 1.3333333333333333
4789.999n 1.0 0.0 1.0 0.3333333333333333 1.3333333333333333
4790n 0.0 0.3333333333333333 0.3333333333333333 0.6666666666666666 0.3333333333333333
4799.999n 0.0 0.3333333333333333 0.3333333333333333 0.6666666666666666 0.3333333333333333
4800n 0.0 0.6666666666666666 0.3333333333333333 0.0 0.5555555555555556
4809.999n 0.0 0.6666666666666666 0.3333333333333333 0.0 0.5555555555555556
4810n 1.0 0.0 0.3333333333333333 1.0 1.1111111111111112
4819.999n 1.0 0.0 0.3333333333333333 1.0 1.1111111111111112
4820n 0.0 0.6666666666666666 0.0 0.0 0.4444444444444444
4829.999n 0.0 0.6666666666666666 0.0 0.0 0.4444444444444444
4830n 0.6666666666666666 0.6666666666666666 0.3333333333333333 0.6666666666666666 1.2222222222222223
4839.999n 0.6666666666666666 0.6666666666666666 0.3333333333333333 0.6666666666666666 1.2222222222222223
4840n 0.6666666666666666 1.0 0.0 0.0 1.3333333333333333
4849.999n 0.6666666666666666 1.0 0.0 0.0 1.3333333333333333
4850n 0.3333333333333333 0.3333333333333333 0.6666666666666666 0.0 0.7777777777777778
4859.999n 0.3333333333333333 0.3333333333333333 0.6666666666666666 0.0 0.7777777777777778
4860n 0.6666666666666666 0.0 0.6666666666666666 0.3333333333333333 0.8888888888888888
4869.999n 0.6666666666666666 0.0 0.6666666666666666 0.3333333333333333 0.8888888888888888
4870n 1.0 0.6666666666666666 0.0 0.3333333333333333 1.4444444444444444
4879.999n 1.0 0.6666666666666666 0.0 0.3333333333333333 1.4444444444444444
4880n 0.6666666666666666 1.0 1.0 0.6666666666666666 1.6666666666666667
4889.999n 0.6666666666666666 1.0 1.0 0.6666666666666666 1.6666666666666667
4890n 0.3333333333333333 0.3333333333333333 1.0 0.6666666666666666 0.8888888888888888
4899.999n 0.3333333333333333 0.3333333333333333 1.0 0.6666666666666666 0.8888888888888888
4900n 1.0 1.0 0.3333333333333333 1.0 1.7777777777777777
4909.999n 1.0 1.0 0.3333333333333333 1.0 1.7777777777777777
4910n 0.6666666666666666 0.6666666666666666 0.3333333333333333 1.0 1.2222222222222223
4919.999n 0.6666666666666666 0.6666666666666666 0.3333333333333333 1.0 1.2222222222222223
4920n 0.6666666666666666 0.3333333333333333 1.0 0.3333333333333333 1.2222222222222223
4929.999n 0.6666666666666666 0.3333333333333333 1.0 0.3333333333333333 1.2222222222222223
4930n 0.0 0.0 0.3333333333333333 0.3333333333333333 0.1111111111111111
4939.999n 0.0 0.0 0.3333333333333333 0.3333333333333333 0.1111111111111111
4940n 0.6666666666666666 1.0 0.0 1.0 1.3333333333333333
4949.999n 0.6666666666666666 1.0 0.0 1.0 1.3333333333333333
4950n 0.6666666666666666 0.0 0.0 0.0 0.6666666666666666
4959.999n 0.6666666666666666 0.0 0.0 0.0 0.6666666666666666
4960n 0.6666666666666666 0.0 1.0 1.0 1.0
4969.999n 0.6666666666666666 0.0 1.0 1.0 1.0
4970n 0.6666666666666666 1.0 0.3333333333333333 0.0 1.4444444444444444
4979.999n 0.6666666666666666 1.0 0.3333333333333333 0.0 1.4444444444444444
4980n 1.0 0.3333333333333333 0.6666666666666666 0.6666666666666666 1.4444444444444444
4989.999n 1.0 0.3333333333333333 0.6666666666666666 0.6666666666666666 1.4444444444444444
4990n 1.0 0.6666666666666666 0.6666666666666666 1.0 1.6666666666666667
4999.999n 1.0 0.6666666666666666 0.6666666666666666 1.0 1.6666666666666667
5000n 1.0 1.0 0.3333333333333333 1.0 1.7777777777777777
5009.999n 1.0 1.0 0.3333333333333333 1.0 1.7777777777777777
5010n 0.0 0.0 0.3333333333333333 0.6666666666666666 0.1111111111111111
5019.999n 0.0 0.0 0.3333333333333333 0.6666666666666666 0.1111111111111111
5020n 0.0 0.6666666666666666 1.0 0.0 0.7777777777777778
5029.999n 0.0 0.6666666666666666 1.0 0.0 0.7777777777777778
5030n 0.3333333333333333 0.0 1.0 0.3333333333333333 0.6666666666666666
5039.999n 0.3333333333333333 0.0 1.0 0.3333333333333333 0.6666666666666666
5040n 0.0 0.0 0.6666666666666666 0.0 0.2222222222222222
5049.999n 0.0 0.0 0.6666666666666666 0.0 0.2222222222222222
5050n 1.0 0.0 0.3333333333333333 1.0 1.1111111111111112
5059.999n 1.0 0.0 0.3333333333333333 1.0 1.1111111111111112
5060n 1.0 1.0 1.0 0.0 2.0
5069.999n 1.0 1.0 1.0 0.0 2.0
5070n 1.0 0.6666666666666666 0.6666666666666666 0.3333333333333333 1.6666666666666667
5079.999n 1.0 0.6666666666666666 0.6666666666666666 0.3333333333333333 1.6666666666666667
5080n 0.3333333333333333 0.0 0.0 0.6666666666666666 0.3333333333333333
5089.999n 0.3333333333333333 0.0 0.0 0.6666666666666666 0.3333333333333333
5090n 1.0 0.3333333333333333 1.0 0.0 1.5555555555555556
5099.999n 1.0 0.3333333333333333 1.0 0.0 1.5555555555555556
5100n 1.0 0.0 0.3333333333333333 0.6666666666666666 1.1111111111111112
5109.999n 1.0 0.0 0.3333333333333333 0.6666666666666666 1.1111111111111112
5110n 0.6666666666666666 0.3333333333333333 1.0 1.0 1.2222222222222223
5119.999n 0.6666666666666666 0.3333333333333333 1.0 1.0 1.2222222222222223
5120n 1.0 0.6666666666666666 0.6666666666666666 0.3333333333333333 1.6666666666666667
5129.999n 1.0 0.6666666666666666 0.6666666666666666 0.3333333333333333 1.6666666666666667
5130n 0.6666666666666666 0.3333333333333333 0.3333333333333333 0.6666666666666666 1.0
5139.999n 0.6666666666666666 0.3333333333333333 0.3333333333333333 0.6666666666666666 1.0
5140n 0.0 0.3333333333333333 0.0 0.0 0.2222222222222222
5149.999n 0.0 0.3333333333333333 0.0 0.0 0.2222222222222222
5150n 0.3333333333333333 1.0 0.0 0.3333333333333333 1.0
5159.999n 0.3333333333333333 1.0 0.0 0.3333333333333333 1.0
5160n 0.0 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.5555555555555556
5169.999n 0.0 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.5555555555555556
5170n 0.3333333333333333 0.0 0.0 0.0 0.3333333333333333
5179.999n 0.3333333333333333 0.0 0.0 0.0 0.3333333333333333
5180n 0.0 0.3333333333333333 0.6666666666666666 1.0 0.4444444444444444
5189.999n 0.0 0.3333333333333333 0.6666666666666666 1.0 0.4444444444444444
5190n 0.6666666666666666 0.6666666666666666 0.6666666666666666 0.0 1.3333333333333333
5199.999n 0.6666666666666666 0.6666666666666666 0.6666666666666666 0.0 1.3333333333333333
5200n 0.6666666666666666 0.0 0.6666666666666666 0.0 0.8888888888888888
5209.999n 0.6666666666666666 0.0 0.6666666666666666 0.0 0.8888888888888888
5210n 0.6666666666666666 1.0 0.0 0.6666666666666666 1.3333333333333333
5219.999n 0.6666666666666666 1.0 0.0 0.6666666666666666 1.3333333333333333
5220n 0.6666666666666666 0.6666666666666666 0.3333333333333333 0.6666666666666666 1.2222222222222223
5229.999n 0.6666666666666666 0.6666666666666666 0.3333333333333333 0.6666666666666666 1.2222222222222223
5230n 0.6666666666666666 0.6666666666666666 0.0 0.6666666666666666 1.1111111111111112
5239.999n 0.6666666666666666 0.6666666666666666 0.0 0.6666666666666666 1.1111111111111112
5240n 0.0 1.0 0.3333333333333333 0.6666666666666666 0.7777777777777778
5249.999n 0.0 1.0 0.3333333333333333 0.6666666666666666 0.7777777777777778
5250n 0.6666666666666666 0.6666666666666666 0.6666666666666666 0.0 1.3333333333333333
5259.999n 0.6666666666666666 0.6666666666666666 0.6666666666666666 0.0 1.3333333333333333
5260n 0.0 0.6666666666666666 0.0 0.3333333333333333 0.4444444444444444
5269.999n 0.0 0.6666666666666666 0.0 0.3333333333333333 0.4444444444444444
5270n 0.0 1.0 0.6666666666666666 1.0 0.8888888888888888
5279.999n 0.0 1.0 0.6666666666666666 1.0 0.8888888888888888
5280n 0.3333333333333333 0.6666666666666666 1.0 0.0 1.1111111111111112
5289.999n 0.3333333333333333 0.6666666666666666 1.0 0.0 1.1111111111111112
5290n 0.3333333333333333 0.0 0.3333333333333333 1.0 0.4444444444444444
5299.999n 0.3333333333333333 0.0 0.3333333333333333 1.0 0.4444444444444444
5300n 1.0 0.3333333333333333 0.3333333333333333 0.6666666666666666 1.3333333333333333
5309.999n 1.0 0.3333333333333333 0.3333333333333333 0.6666666666666666 1.3333333333333333
5310n 1.0 0.0 0.3333333333333333 0.6666666666666666 1.1111111111111112
5319.999n 1.0 0.0 0.3333333333333333 0.6666666666666666 1.1111111111111112
5320n 0.6666666666666666 0.6666666666666666 0.3333333333333333 0.3333333333333333 1.2222222222222223
5329.999n 0.6666666666666666 0.6666666666666666 0.3333333333333333 0.3333333333333333 1.2222222222222223
5330n 0.3333333333333333 1.0 1.0 0.0 1.3333333333333333
5339.999n 0.3333333333333333 1.0 1.0 0.0 1.3333333333333333
5340n 0.6666666666666666 0.3333333333333333 0.3333333333333333 0.3333333333333333 1.0
5349.999n 0.6666666666666666 0.3333333333333333 0.3333333333333333 0.3333333333333333 1.0
5350n 0.0 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.5555555555555556
5359.999n 0.0 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.5555555555555556
5360n 0.6666666666666666 0.3333333333333333 0.6666666666666666 1.0 1.1111111111111112
5369.999n 0.6666666666666666 0.3333333333333333 0.6666666666666666 1.0 1.1111111111111112
5370n 0.6666666666666666 0.3333333333333333 1.0 0.0 1.2222222222222223
5379.999n 0.6666666666666666 0.3333333333333333 1.0 0.0 1.2222222222222223
5380n 0.0 0.0 0.6666666666666666 0.6666666666666666 0.2222222222222222
5389.999n 0.0 0.0 0.6666666666666666 0.6666666666666666 0.2222222222222222
5390n 1.0 0.6666666666666666 0.6666666666666666 0.3333333333333333 1.6666666666666667
5399.999n 1.0 0.6666666666666666 0.6666666666666666 0.3333333333333333 1.6666666666666667
5400n 0.3333333333333333 1.0 0.6666666666666666 1.0 1.2222222222222223
5409.999n 0.3333333333333333 1.0 0.6666666666666666 1.0 1.2222222222222223
5410n 0.0 0.6666666666666666 0.6666666666666666 0.6666666666666666 0.6666666666666666
5419.999n 0.0 0.6666666666666666 0.6666666666666666 0.6666666666666666 0.6666666666666666
5420n 1.0 0.6666666666666666 0.3333333333333333 0.3333333333333333 1.5555555555555556
5429.999n 1.0 0.6666666666666666 0.3333333333333333 0.3333333333333333 1.5555555555555556
5430n 0.6666666666666666 0.3333333333333333 0.0 0.3333333333333333 0.8888888888888888
5439.999n 0.6666666666666666 0.3333333333333333 0.0 0.3333333333333333 0.8888888888888888
5440n 0.3333333333333333 1.0 0.0 0.0 1.0
5449.999n 0.3333333333333333 1.0 0.0 0.0 1.0
5450n 1.0 1.0 0.3333333333333333 0.3333333333333333 1.7777777777777777
5459.999n 1.0 1.0 0.3333333333333333 0.3333333333333333 1.7777777777777777
5460n 0.6666666666666666 0.6666666666666666 1.0 0.0 1.4444444444444444
5469.999n 0.6666666666666666 0.6666666666666666 1.0 0.0 1.4444444444444444
5470n 1.0 0.0 0.3333333333333333 0.0 1.1111111111111112
5479.999n 1.0 0.0 0.3333333333333333 0.0 1.1111111111111112
5480n 0.0 0.6666666666666666 0.0 0.3333333333333333 0.4444444444444444
5489.999n 0.0 0.6666666666666666 0.0 0.3333333333333333 0.4444444444444444
5490n 0.6666666666666666 0.0 1.0 0.3333333333333333 1.0
5499.999n 0.6666666666666666 0.0 1.0 0.3333333333333333 1.0
5500n 0.6666666666666666 0.0 0.3333333333333333 0.6666666666666666 0.7777777777777778
5509.999n 0.6666666666666666 0.0 0.3333333333333333 0.6666666666666666 0.7777777777777778
5510n 0.6666666666666666 1.0 1.0 1.0 1.6666666666666667
5519.999n 0.6666666666666666 1.0 1.0 1.0 1.6666666666666667
5520n 0.3333333333333333 0.0 0.6666666666666666 0.3333333333333333 0.5555555555555556
5529.999n 0.3333333333333333 0.0 0.6666666666666666 0.3333333333333333 0.5555555555555556
5530n 0.6666666666666666 0.0 0.3333333333333333 1.0 0.7777777777777778
5539.999n 0.6666666666666666 0.0 0.3333333333333333 1.0 0.7777777777777778
5540n 0.6666666666666666 0.0 0.6666666666666666 0.0 0.8888888888888888
5549.999n 0.6666666666666666 0.0 0.6666666666666666 0.0 0.8888888888888888
5550n 0.0 0.6666666666666666 0.6666666666666666 0.0 0.6666666666666666
5559.999n 0.0 0.6666666666666666 0.6666666666666666 0.0 0.6666666666666666
5560n 1.0 0.6666666666666666 0.0 0.6666666666666666 1.4444444444444444
5569.999n 1.0 0.6666666666666666 0.0 0.6666666666666666 1.4444444444444444
5570n 0.0 1.0 0.3333333333333333 0.3333333333333333 0.7777777777777778
5579.999n 0.0 1.0 0.3333333333333333 0.3333333333333333 0.7777777777777778
5580n 0.0 0.0 0.3333333333333333 0.0 0.1111111111111111
5589.999n 0.0 0.0 0.3333333333333333 0.0 0.1111111111111111
5590n 0.3333333333333333 0.3333333333333333 0.3333333333333333 1.0 0.6666666666666666
5599.999n 0.3333333333333333 0.3333333333333333 0.3333333333333333 1.0 0.6666666666666666
5600n 0.6666666666666666 0.3333333333333333 0.0 0.6666666666666666 0.8888888888888888
5609.999n 0.6666666666666666 0.3333333333333333 0.0 0.6666666666666666 0.8888888888888888
5610n 0.3333333333333333 1.0 1.0 0.0 1.3333333333333333
5619.999n 0.3333333333333333 1.0 1.0 0.0 1.3333333333333333
5620n 0.0 1.0 0.3333333333333333 0.3333333333333333 0.7777777777777778
5629.999n 0.0 1.0 0.3333333333333333 0.3333333333333333 0.7777777777777778
5630n 0.3333333333333333 1.0 0.6666666666666666 0.0 1.2222222222222223
5639.999n 0.3333333333333333 1.0 0.6666666666666666 0.0 1.2222222222222223
5640n 0.0 0.0 0.6666666666666666 0.3333333333333333 0.2222222222222222
5649.999n 0.0 0.0 0.6666666666666666 0.3333333333333333 0.2222222222222222
5650n 0.6666666666666666 0.6666666666666666 0.6666666666666666 0.3333333333333333 1.3333333333333333
5659.999n 0.6666666666666666 0.6666666666666666 0.6666666666666666 0.3333333333333333 1.3333333333333333
5660n 0.6666666666666666 0.3333333333333333 0.3333333333333333 0.3333333333333333 1.0
5669.999n 0.6666666666666666 0.3333333333333333 0.3333333333333333 0.3333333333333333 1.0
5670n 0.3333333333333333 1.0 1.0 0.0 1.3333333333333333
5679.999n 0.3333333333333333 1.0 1.0 0.0 1.3333333333333333
5680n 0.0 0.3333333333333333 1.0 0.3333333333333333 0.5555555555555556
5689.999n 0.0 0.3333333333333333 1.0 0.3333333333333333 0.5555555555555556
5690n 1.0 1.0 0.3333333333333333 0.3333333333333333 1.7777777777777777
5699.999n 1.0 1.0 0.3333333333333333 0.3333333333333333 1.7777777777777777
5700n 1.0 0.3333333333333333 0.6666666666666666 0.0 1.4444444444444444
5709.999n 1.0 0.3333333333333333 0.6666666666666666 0.0 1.4444444444444444
5710n 0.6666666666666666 0.6666666666666666 1.0 0.6666666666666666 1.4444444444444444
5719.999n 0.6666666666666666 0.6666666666666666 1.0 0.6666666666666666 1.4444444444444444
5720n 0.6666666666666666 0.3333333333333333 1.0 0.6666666666666666 1.2222222222222223
5729.999n 0.6666666666666666 0.3333333333333333 1.0 0.6666666666666666 1.2222222222222223
5730n 0.3333333333333333 0.0 0.0 0.6666666666666666 0.3333333333333333
5739.999n 0.3333333333333333 0.0 0.0 0.6666666666666666 0.3333333333333333
5740n 0.6666666666666666 0.6666666666666666 0.6666666666666666 1.0 1.3333333333333333
5749.999n 0.6666666666666666 0.6666666666666666 0.6666666666666666 1.0 1.3333333333333333
5750n 1.0 0.0 0.6666666666666666 1.0 1.2222222222222223
5759.999n 1.0 0.0 0.6666666666666666 1.0 1.2222222222222223
5760n 1.0 0.0 0.6666666666666666 0.0 1.2222222222222223
5769.999n 1.0 0.0 0.6666666666666666 0.0 1.2222222222222223
5770n 1.0 1.0 0.0 0.0 1.6666666666666667
5779.999n 1.0 1.0 0.0 0.0 1.6666666666666667
5780n 0.6666666666666666 0.6666666666666666 0.3333333333333333 0.3333333333333333 1.2222222222222223
5789.999n 0.6666666666666666 0.6666666666666666 0.3333333333333333 0.3333333333333333 1.2222222222222223
5790n 0.6666666666666666 0.0 1.0 0.3333333333333333 1.0
5799.999n 0.6666666666666666 0.0 1.0 0.3333333333333333 1.0
5800n 0.3333333333333333 0.0 0.0 0.0 0.3333333333333333
5809.999n 0.3333333333333333 0.0 0.0 0.0 0.3333333333333333
5810n 0.0 0.0 0.3333333333333333 0.3333333333333333 0.1111111111111111
5819.999n 0.0 0.0 0.3333333333333333 0.3333333333333333 0.1111111111111111
5820n 0.6666666666666666 1.0 1.0 0.3333333333333333 1.6666666666666667
5829.999n 0.6666666666666666 1.0 1.0 0.3333333333333333 1.6666666666666667
5830n 0.0 1.0 1.0 0.6666666666666666 1.0
5839.999n 0.0 1.0 1.0 0.6666666666666666 1.0
5840n 0.6666666666666666 0.6666666666666666 0.3333333333333333 0.0 1.2222222222222223
5849.999n 0.6666666666666666 0.6666666666666666 0.3333333333333333 0.0 1.2222222222222223
5850n 0.3333333333333333 1.0 0.6666666666666666 0.6666666666666666 1.2222222222222223
5859.999n 0.3333333333333333 1.0 0.6666666666666666 0.6666666666666666 1.2222222222222223
5860n 0.6666666666666666 0.3333333333333333 0.0 0.6666666666666666 0.8888888888888888
5869.999n 0.6666666666666666 0.3333333333333333 0.0 0.6666666666666666 0.8888888888888888
5870n 0.3333333333333333 0.0 0.6666666666666666 0.3333333333333333 0.5555555555555556
5879.999n 0.3333333333333333 0.0 0.6666666666666666 0.3333333333333333 0.5555555555555556
5880n 0.3333333333333333 0.3333333333333333 1.0 0.6666666666666666 0.8888888888888888
5889.999n 0.3333333333333333 0.3333333333333333 1.0 0.6666666666666666 0.8888888888888888
5890n 1.0 0.0 0.0 0.3333333333333333 1.0
5899.999n 1.0 0.0 0.0 0.3333333333333333 1.0
5900n 1.0 0.6666666666666666 1.0 0.3333333333333333 1.7777777777777777
5909.999n 1.0 0.6666666666666666 1.0 0.3333333333333333 1.7777777777777777
5910n 0.6666666666666666 0.0 0.6666666666666666 1.0 0.8888888888888888
5919.999n 0.6666666666666666 0.0 0.6666666666666666 1.0 0.8888888888888888
5920n 0.6666666666666666 0.0 0.0 0.3333333333333333 0.6666666666666666
5929.999n 0.6666666666666666 0.0 0.0 0.3333333333333333 0.6666666666666666
5930n 0.3333333333333333 0.3333333333333333 1.0 1.0 0.8888888888888888
5939.999n 0.3333333333333333 0.3333333333333333 1.0 1.0 0.8888888888888888
5940n 0.0 1.0 1.0 1.0 1.0
5949.999n 0.0 1.0 1.0 1.0 1.0
5950n 0.6666666666666666 1.0 0.3333333333333333 0.3333333333333333 1.4444444444444444
5959.999n 0.6666666666666666 1.0 0.3333333333333333 0.3333333333333333 1.4444444444444444
5960n 0.0 0.0 0.3333333333333333 0.0 0.1111111111111111
5969.999n 0.0 0.0 0.3333333333333333 0.0 0.1111111111111111
5970n 0.6666666666666666 0.6666666666666666 0.0 0.0 1.1111111111111112
5979.999n 0.6666666666666666 0.6666666666666666 0.0 0.0 1.1111111111111112
5980n 0.0 0.6666666666666666 0.0 0.6666666666666666 0.4444444444444444
5989.999n 0.0 0.6666666666666666 0.0 0.6666666666666666 0.4444444444444444
5990n 0.0 0.3333333333333333 0.6666666666666666 1.0 0.4444444444444444
5999.999n 0.0 0.3333333333333333 0.6666666666666666 1.0 0.4444444444444444
6000n 1.0 0.0 1.0 1.0 1.3333333333333333
6009.999n 1.0 0.0 1.0 1.0 1.3333333333333333
6010n 1.0 1.0 0.3333333333333333 0.6666666666666666 1.7777777777777777
6019.999n 1.0 1.0 0.3333333333333333 0.6666666666666666 1.7777777777777777
6020n 0.6666666666666666 0.6666666666666666 0.0 1.0 1.1111111111111112
6029.999n 0.6666666666666666 0.6666666666666666 0.0 1.0 1.1111111111111112
6030n 0.0 0.6666666666666666 0.0 0.6666666666666666 0.4444444444444444
6039.999n 0.0 0.6666666666666666 0.0 0.6666666666666666 0.4444444444444444
6040n 0.3333333333333333 0.6666666666666666 0.3333333333333333 1.0 0.8888888888888888
6049.999n 0.3333333333333333 0.6666666666666666 0.3333333333333333 1.0 0.8888888888888888
6050n 1.0 0.3333333333333333 0.0 0.3333333333333333 1.2222222222222223
6059.999n 1.0 0.3333333333333333 0.0 0.3333333333333333 1.2222222222222223
6060n 1.0 0.3333333333333333 0.3333333333333333 0.0 1.3333333333333333
6069.999n 1.0 0.3333333333333333 0.3333333333333333 0.0 1.3333333333333333
6070n 0.6666666666666666 0.3333333333333333 0.0 0.6666666666666666 0.8888888888888888
6079.999n 0.6666666666666666 0.3333333333333333 0.0 0.6666666666666666 0.8888888888888888
6080n 1.0 0.0 0.6666666666666666 0.0 1.2222222222222223
6089.999n 1.0 0.0 0.6666666666666666 0.0 1.2222222222222223
6090n 0.3333333333333333 0.0 0.0 0.3333333333333333 0.3333333333333333
6099.999n 0.3333333333333333 0.0 0.0 0.3333333333333333 0.3333333333333333
6100n 1.0 1.0 0.6666666666666666 0.6666666666666666 1.8888888888888888
6109.999n 1.0 1.0 0.6666666666666666 0.6666666666666666 1.8888888888888888
6110n 0.3333333333333333 0.3333333333333333 1.0 0.6666666666666666 0.8888888888888888
6119.999n 0.3333333333333333 0.3333333333333333 1.0 0.6666666666666666 0.8888888888888888
6120n 0.0 0.0 0.0 0.0 0.0
6129.999n 0.0 0.0 0.0 0.0 0.0
6130n 1.0 0.6666666666666666 0.0 0.3333333333333333 1.4444444444444444
6139.999n 1.0 0.6666666666666666 0.0 0.3333333333333333 1.4444444444444444
6140n 0.3333333333333333 1.0 0.0 1.0 1.0
6149.999n 0.3333333333333333 1.0 0.0 1.0 1.0
6150n 0.0 0.0 0.3333333333333333 0.6666666666666666 0.1111111111111111
6159.999n 0.0 0.0 0.3333333333333333 0.6666666666666666 0.1111111111111111
6160n 1.0 0.3333333333333333 0.6666666666666666 0.3333333333333333 1.4444444444444444
6169.999n 1.0 0.3333333333333333 0.6666666666666666 0.3333333333333333 1.4444444444444444
6170n 0.6666666666666666 1.0 0.3333333333333333 0.6666666666666666 1.4444444444444444
6179.999n 0.6666666666666666 1.0 0.3333333333333333 0.6666666666666666 1.4444444444444444
6180n 0.3333333333333333 0.6666666666666666 0.6666666666666666 1.0 1.0
6189.999n 0.3333333333333333 0.6666666666666666 0.6666666666666666 1.0 1.0
6190n 0.0 0.3333333333333333 1.0 1.0 0.5555555555555556
6199.999n 0.0 0.3333333333333333 1.0 1.0 0.5555555555555556
6200n 1.0 0.6666666666666666 1.0 1.0 1.7777777777777777
6209.999n 1.0 0.6666666666666666 1.0 1.0 1.7777777777777777
6210n 0.3333333333333333 0.0 0.0 0.3333333333333333 0.3333333333333333
6219.999n 0.3333333333333333 0.0 0.0 0.3333333333333333 0.3333333333333333
6220n 0.0 0.6666666666666666 0.0 0.0 0.4444444444444444
6229.999n 0.0 0.6666666666666666 0.0 0.0 0.4444444444444444
6230n 0.3333333333333333 1.0 0.3333333333333333 0.3333333333333333 1.1111111111111112
6239.999n 0.3333333333333333 1.0 0.3333333333333333 0.3333333333333333 1.1111111111111112
6240n 0.0 0.6666666666666666 0.0 0.3333333333333333 0.4444444444444444
6249.999n 0.0 0.6666666666666666 0.0 0.3333333333333333 0.4444444444444444
6250n 0.0 0.3333333333333333 1.0 0.3333333333333333 0.5555555555555556
6259.999n 0.0 0.3333333333333333 1.0 0.3333333333333333 0.5555555555555556
6260n 0.6666666666666666 0.3333333333333333 0.3333333333333333 0.3333333333333333 1.0
6269.999n 0.6666666666666666 0.3333333333333333 0.3333333333333333 0.3333333333333333 1.0
6270n 0.6666666666666666 0.0 1.0 0.0 1.0
6279.999n 0.6666666666666666 0.0 1.0 0.0 1.0
6280n 1.0 0.6666666666666666 0.6666666666666666 0.0 1.6666666666666667
6289.999n 1.0 0.6666666666666666 0.6666666666666666 0.0 1.6666666666666667
6290n 0.6666666666666666 1.0 1.0 1.0 1.6666666666666667
6299.999n 0.6666666666666666 1.0 1.0 1.0 1.6666666666666667
6300n 0.0 0.3333333333333333 0.0 0.6666666666666666 0.2222222222222222
6309.999n 0.0 0.3333333333333333 0.0 0.6666666666666666 0.2222222222222222
6310n 0.6666666666666666 0.0 1.0 0.0 1.0
6319.999n 0.6666666666666666 0.0 1.0 0.0 1.0
6320n 0.6666666666666666 1.0 0.3333333333333333 1.0 1.4444444444444444
6329.999n 0.6666666666666666 1.0 0.3333333333333333 1.0 1.4444444444444444
6330n 0.3333333333333333 1.0 0.6666666666666666 0.6666666666666666 1.2222222222222223
6339.999n 0.3333333333333333 1.0 0.6666666666666666 0.6666666666666666 1.2222222222222223
6340n 0.6666666666666666 0.6666666666666666 0.6666666666666666 0.6666666666666666 1.3333333333333333
6349.999n 0.6666666666666666 0.6666666666666666 0.6666666666666666 0.6666666666666666 1.3333333333333333
6350n 0.0 0.3333333333333333 0.3333333333333333 0.3333333333333333 0.3333333333333333
6359.999n 0.0 0.3333333333333333 0.3333333333333333 0.3333333333333333 0.3333333333333333
6360n 0.0 1.0 0.3333333333333333 1.0 0.7777777777777778
6369.999n 0.0 1.0 0.3333333333333333 1.0 0.7777777777777778
6370n 0.0 1.0 0.6666666666666666 0.3333333333333333 0.8888888888888888
6379.999n 0.0 1.0 0.6666666666666666 0.3333333333333333 0.8888888888888888
6380n 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.3333333333333333 1.1111111111111112
6389.999n 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.3333333333333333 1.1111111111111112
6390n 1.0 0.3333333333333333 0.0 0.3333333333333333 1.2222222222222223
6399.999n 1.0 0.3333333333333333 0.0 0.3333333333333333 1.2222222222222223
6400n 0.6666666666666666 0.0 0.6666666666666666 1.0 0.8888888888888888
6409.999n 0.6666666666666666 0.0 0.6666666666666666 1.0 0.8888888888888888
6410n 0.0 0.3333333333333333 0.3333333333333333 0.0 0.3333333333333333
6419.999n 0.0 0.3333333333333333 0.3333333333333333 0.0 0.3333333333333333
6420n 0.6666666666666666 1.0 1.0 0.0 1.6666666666666667
6429.999n 0.6666666666666666 1.0 1.0 0.0 1.6666666666666667
6430n 0.6666666666666666 1.0 0.6666666666666666 0.3333333333333333 1.5555555555555556
6439.999n 0.6666666666666666 1.0 0.6666666666666666 0.3333333333333333 1.5555555555555556
6440n 0.6666666666666666 1.0 1.0 0.0 1.6666666666666667
6449.999n 0.6666666666666666 1.0 1.0 0.0 1.6666666666666667
6450n 0.0 0.0 0.6666666666666666 1.0 0.2222222222222222
6459.999n 0.0 0.0 0.6666666666666666 1.0 0.2222222222222222
6460n 0.6666666666666666 0.0 0.0 1.0 0.6666666666666666
6469.999n 0.6666666666666666 0.0 0.0 1.0 0.6666666666666666
6470n 1.0 0.0 1.0 0.3333333333333333 1.3333333333333333
6479.999n 1.0 0.0 1.0 0.3333333333333333 1.3333333333333333
6480n 0.0 1.0 1.0 0.0 1.0
6489.999n 0.0 1.0 1.0 0.0 1.0
6490n 0.0 0.0 0.3333333333333333 1.0 0.1111111111111111
6499.999n 0.0 0.0 0.3333333333333333 1.0 0.1111111111111111
6500n 0.3333333333333333 0.0 0.0 0.3333333333333333 0.3333333333333333
6509.999n 0.3333333333333333 0.0 0.0 0.3333333333333333 0.3333333333333333
6510n 1.0 0.0 0.0 0.0 1.0
6519.999n 1.0 0.0 0.0 0.0 1.0
6520n 0.3333333333333333 1.0 0.0 0.0 1.0
6529.999n 0.3333333333333333 1.0 0.0 0.0 1.0
6530n 1.0 0.6666666666666666 0.3333333333333333 0.3333333333333333 1.5555555555555556
6539.999n 1.0 0.6666666666666666 0.3333333333333333 0.3333333333333333 1.5555555555555556
6540n 0.6666666666666666 0.0 1.0 0.0 1.0
6549.999n 0.6666666666666666 0.0 1.0 0.0 1.0
6550n 0.3333333333333333 0.6666666666666666 0.0 0.3333333333333333 0.7777777777777778
6559.999n 0.3333333333333333 0.6666666666666666 0.0 0.3333333333333333 0.7777777777777778
6560n 0.3333333333333333 0.0 0.6666666666666666 0.3333333333333333 0.5555555555555556
6569.999n 0.3333333333333333 0.0 0.6666666666666666 0.3333333333333333 0.5555555555555556
6570n 0.6666666666666666 1.0 0.6666666666666666 1.0 1.5555555555555556
6579.999n 0.6666666666666666 1.0 0.6666666666666666 1.0 1.5555555555555556
6580n 1.0 0.3333333333333333 0.3333333333333333 0.3333333333333333 1.3333333333333333
6589.999n 1.0 0.3333333333333333 0.3333333333333333 0.3333333333333333 1.3333333333333333
6590n 1.0 0.3333333333333333 1.0 0.0 1.5555555555555556
6599.999n 1.0 0.3333333333333333 1.0 0.0 1.5555555555555556
6600n 0.3333333333333333 0.3333333333333333 0.0 0.0 0.5555555555555556
6609.999n 0.3333333333333333 0.3333333333333333 0.0 0.0 0.5555555555555556
6610n 1.0 0.3333333333333333 0.6666666666666666 0.0 1.4444444444444444
6619.999n 1.0 0.3333333333333333 0.6666666666666666 0.0 1.4444444444444444
6620n 0.0 0.0 0.0 0.6666666666666666 0.0
6629.999n 0.0 0.0 0.0 0.6666666666666666 0.0
6630n 0.6666666666666666 0.0 0.6666666666666666 0.6666666666666666 0.8888888888888888
6639.999n 0.6666666666666666 0.0 0.6666666666666666 0.6666666666666666 0.8888888888888888
6640n 1.0 1.0 0.3333333333333333 0.6666666666666666 1.7777777777777777
6649.999n 1.0 1.0 0.3333333333333333 0.6666666666666666 1.7777777777777777
6650n 0.6666666666666666 0.6666666666666666 1.0 0.6666666666666666 1.4444444444444444
6659.999n 0.6666666666666666 0.6666666666666666 1.0 0.6666666666666666 1.4444444444444444
6660n 0.0 1.0 0.0 1.0 0.6666666666666666
6669.999n 0.0 1.0 0.0 1.0 0.6666666666666666
6670n 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.6666666666666666 1.1111111111111112
6679.999n 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.6666666666666666 1.1111111111111112
6680n 1.0 0.3333333333333333 0.6666666666666666 0.0 1.4444444444444444
6689.999n 1.0 0.3333333333333333 0.6666666666666666 0.0 1.4444444444444444
6690n 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.6666666666666666 1.1111111111111112
6699.999n 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.6666666666666666 1.1111111111111112
6700n 0.0 0.3333333333333333 0.0 0.3333333333333333 0.2222222222222222
6709.999n 0.0 0.3333333333333333 0.0 0.3333333333333333 0.2222222222222222
6710n 0.3333333333333333 0.6666666666666666 0.0 0.6666666666666666 0.7777777777777778
6719.999n 0.3333333333333333 0.6666666666666666 0.0 0.6666666666666666 0.7777777777777778
6720n 1.0 0.3333333333333333 0.0 0.3333333333333333 1.2222222222222223
6729.999n 1.0 0.3333333333333333 0.0 0.3333333333333333 1.2222222222222223
6730n 0.3333333333333333 0.6666666666666666 0.3333333333333333 0.3333333333333333 0.8888888888888888
6739.999n 0.3333333333333333 0.6666666666666666 0.3333333333333333 0.3333333333333333 0.8888888888888888
6740n 0.3333333333333333 0.6666666666666666 0.3333333333333333 1.0 0.8888888888888888
6749.999n 0.3333333333333333 0.6666666666666666 0.3333333333333333 1.0 0.8888888888888888
6750n 0.0 0.6666666666666666 1.0 1.0 0.7777777777777778
6759.999n 0.0 0.6666666666666666 1.0 1.0 0.7777777777777778
6760n 0.0 0.6666666666666666 0.0 0.0 0.4444444444444444
6769.999n 0.0 0.6666666666666666 0.0 0.0 0.4444444444444444
6770n 0.0 0.3333333333333333 0.6666666666666666 0.0 0.4444444444444444
6779.999n 0.0 0.3333333333333333 0.6666666666666666 0.0 0.4444444444444444
6780n 0.3333333333333333 1.0 0.6666666666666666 0.3333333333333333 1.2222222222222223
6789.999n 0.3333333333333333 1.0 0.6666666666666666 0.3333333333333333 1.2222222222222223
6790n 0.6666666666666666 1.0 0.6666666666666666 0.3333333333333333 1.5555555555555556
6799.999n 0.6666666666666666 1.0 0.6666666666666666 0.3333333333333333 1.5555555555555556
6800n 0.6666666666666666 1.0 0.3333333333333333 0.6666666666666666 1.4444444444444444
6809.999n 0.6666666666666666 1.0 0.3333333333333333 0.6666666666666666 1.4444444444444444
6810n 1.0 0.6666666666666666 0.0 0.6666666666666666 1.4444444444444444
6819.999n 1.0 0.6666666666666666 0.0 0.6666666666666666 1.4444444444444444
6820n 1.0 0.0 0.3333333333333333 0.3333333333333333 1.1111111111111112
6829.999n 1.0 0.0 0.3333333333333333 0.3333333333333333 1.1111111111111112
6830n 0.3333333333333333 0.0 0.3333333333333333 0.0 0.4444444444444444
6839.999n 0.3333333333333333 0.0 0.3333333333333333 0.0 0.4444444444444444
6840n 0.0 0.0 0.6666666666666666 0.0 0.2222222222222222
6849.999n 0.0 0.0 0.6666666666666666 0.0 0.2222222222222222
6850n 1.0 0.3333333333333333 0.3333333333333333 0.0 1.3333333333333333
6859.999n 1.0 0.3333333333333333 0.3333333333333333 0.0 1.3333333333333333
6860n 0.0 0.3333333333333333 1.0 1.0 0.5555555555555556
6869.999n 0.0 0.3333333333333333 1.0 1.0 0.5555555555555556
6870n 1.0 0.3333333333333333 0.3333333333333333 1.0 1.3333333333333333
6879.999n 1.0 0.3333333333333333 0.3333333333333333 1.0 1.3333333333333333
6880n 1.0 0.3333333333333333 0.6666666666666666 0.3333333333333333 1.4444444444444444
6889.999n 1.0 0.3333333333333333 0.6666666666666666 0.3333333333333333 1.4444444444444444
6890n 1.0 0.3333333333333333 1.0 0.0 1.5555555555555556
6899.999n 1.0 0.3333333333333333 1.0 0.0 1.5555555555555556
6900n 0.0 0.6666666666666666 0.3333333333333333 0.0 0.5555555555555556
6909.999n 0.0 0.6666666666666666 0.3333333333333333 0.0 0.5555555555555556
6910n 0.6666666666666666 0.6666666666666666 0.0 0.6666666666666666 1.1111111111111112
6919.999n 0.6666666666666666 0.6666666666666666 0.0 0.6666666666666666 1.1111111111111112
6920n 0.0 0.3333333333333333 0.6666666666666666 1.0 0.4444444444444444
6929.999n 0.0 0.3333333333333333 0.6666666666666666 1.0 0.4444444444444444
6930n 0.0 0.3333333333333333 0.0 0.0 0.2222222222222222
6939.999n 0.0 0.3333333333333333 0.0 0.0 0.2222222222222222
6940n 1.0 1.0 0.6666666666666666 1.0 1.8888888888888888
6949.999n 1.0 1.0 0.6666666666666666 1.0 1.8888888888888888
6950n 0.6666666666666666 0.3333333333333333 0.0 0.0 0.8888888888888888
6959.999n 0.6666666666666666 0.3333333333333333 0.0 0.0 0.8888888888888888
6960n 0.0 0.6666666666666666 0.3333333333333333 0.0 0.5555555555555556
6969.999n 0.0 0.6666666666666666 0.3333333333333333 0.0 0.5555555555555556
6970n 1.0 0.3333333333333333 0.6666666666666666 1.0 1.4444444444444444
6979.999n 1.0 0.3333333333333333 0.6666666666666666 1.0 1.4444444444444444
6980n 0.0 0.6666666666666666 1.0 1.0 0.7777777777777778
6989.999n 0.0 0.6666666666666666 1.0 1.0 0.7777777777777778
6990n 0.0 0.3333333333333333 0.3333333333333333 0.6666666666666666 0.3333333333333333
6999.999n 0.0 0.3333333333333333 0.3333333333333333 0.6666666666666666 0.3333333333333333
7000n 1.0 0.0 1.0 0.0 1.3333333333333333
7009.999n 1.0 0.0 1.0 0.0 1.3333333333333333
7010n 0.3333333333333333 0.3333333333333333 1.0 1.0 0.8888888888888888
7019.999n 0.3333333333333333 0.3333333333333333 1.0 1.0 0.8888888888888888
7020n 0.0 0.6666666666666666 1.0 0.3333333333333333 0.7777777777777778
7029.999n 0.0 0.6666666666666666 1.0 0.3333333333333333 0.7777777777777778
7030n 0.6666666666666666 0.0 0.6666666666666666 0.0 0.8888888888888888
7039.999n 0.6666666666666666 0.0 0.6666666666666666 0.0 0.8888888888888888
7040n 1.0 0.0 1.0 0.0 1.3333333333333333
7049.999n 1.0 0.0 1.0 0.0 1.3333333333333333
7050n 1.0 1.0 1.0 0.6666666666666666 2.0
7059.999n 1.0 1.0 1.0 0.6666666666666666 2.0
7060n 0.6666666666666666 1.0 0.6666666666666666 0.6666666666666666 1.5555555555555556
7069.999n 0.6666666666666666 1.0 0.6666666666666666 0.6666666666666666 1.5555555555555556
7070n 0.0 0.3333333333333333 0.3333333333333333 0.6666666666666666 0.3333333333333333
7079.999n 0.0 0.3333333333333333 0.3333333333333333 0.6666666666666666 0.3333333333333333
7080n 0.6666666666666666 1.0 0.6666666666666666 0.0 1.5555555555555556
7089.999n 0.6666666666666666 1.0 0.6666666666666666 0.0 1.5555555555555556
7090n 0.3333333333333333 1.0 0.6666666666666666 1.0 1.2222222222222223
7099.999n 0.3333333333333333 1.0 0.6666666666666666 1.0 1.2222222222222223
7100n 0.0 1.0 0.0 0.0 0.6666666666666666
7109.999n 0.0 1.0 0.0 0.0 0.6666666666666666
7110n 0.6666666666666666 1.0 0.3333333333333333 0.0 1.4444444444444444
7119.999n 0.6666666666666666 1.0 0.3333333333333333 0.0 1.4444444444444444
7120n 0.3333333333333333 0.6666666666666666 1.0 1.0 1.1111111111111112
7129.999n 0.3333333333333333 0.6666666666666666 1.0 1.0 1.1111111111111112
7130n 0.0 0.6666666666666666 0.3333333333333333 1.0 0.5555555555555556
7139.999n 0.0 0.6666666666666666 0.3333333333333333 1.0 0.5555555555555556
7140n 0.3333333333333333 1.0 1.0 0.3333333333333333 1.3333333333333333
7149.999n 0.3333333333333333 1.0 1.0 0.3333333333333333 1.3333333333333333
7150n 1.0 0.3333333333333333 1.0 0.0 1.5555555555555556
7159.999n 1.0 0.3333333333333333 1.0 0.0 1.5555555555555556
7160n 0.3333333333333333 0.6666666666666666 0.0 1.0 0.7777777777777778
7169.999n 0.3333333333333333 0.6666666666666666 0.0 1.0 0.7777777777777778
7170n 0.0 0.3333333333333333 0.3333333333333333 1.0 0.3333333333333333
7179.999n 0.0 0.3333333333333333 0.3333333333333333 1.0 0.3333333333333333
7180n 0.0 1.0 0.3333333333333333 1.0 0.7777777777777778
7189.999n 0.0 1.0 0.3333333333333333 1.0 0.7777777777777778
7190n 0.3333333333333333 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.8888888888888888
7199.999n 0.3333333333333333 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.8888888888888888
7200n 0.0 1.0 0.6666666666666666 1.0 0.8888888888888888
7209.999n 0.0 1.0 0.6666666666666666 1.0 0.8888888888888888
7210n 1.0 0.3333333333333333 0.3333333333333333 0.3333333333333333 1.3333333333333333
7219.999n 1.0 0.3333333333333333 0.3333333333333333 0.3333333333333333 1.3333333333333333
7220n 0.0 0.6666666666666666 1.0 1.0 0.7777777777777778
7229.999n 0.0 0.6666666666666666 1.0 1.0 0.7777777777777778
7230n 0.6666666666666666 0.6666666666666666 0.0 0.6666666666666666 1.1111111111111112
7239.999n 0.6666666666666666 0.6666666666666666 0.0 0.6666666666666666 1.1111111111111112
7240n 1.0 0.0 0.3333333333333333 1.0 1.1111111111111112
7249.999n 1.0 0.0 0.3333333333333333 1.0 1.1111111111111112
7250n 0.6666666666666666 0.6666666666666666 0.6666666666666666 0.3333333333333333 1.3333333333333333
7259.999n 0.6666666666666666 0.6666666666666666 0.6666666666666666 0.3333333333333333 1.3333333333333333
7260n 0.0 1.0 0.6666666666666666 0.0 0.8888888888888888
7269.999n 0.0 1.0 0.6666666666666666 0.0 0.8888888888888888
7270n 0.6666666666666666 0.0 1.0 0.6666666666666666 1.0
7279.999n 0.6666666666666666 0.0 1.0 0.6666666666666666 1.0
7280n 0.0 0.3333333333333333 0.0 0.3333333333333333 0.2222222222222222
7289.999n 0.0 0.3333333333333333 0.0 0.3333333333333333 0.2222222222222222
7290n 0.0 0.0 0.3333333333333333 1.0 0.1111111111111111
7299.999n 0.0 0.0 0.3333333333333333 1.0 0.1111111111111111
7300n 0.3333333333333333 0.0 0.6666666666666666 0.6666666666666666 0.5555555555555556
7309.999n 0.3333333333333333 0.0 0.6666666666666666 0.6666666666666666 0.5555555555555556
7310n 1.0 0.6666666666666666 0.0 0.0 1.4444444444444444
7319.999n 1.0 0.6666666666666666 0.0 0.0 1.4444444444444444
7320n 0.3333333333333333 0.6666666666666666 0.0 0.0 0.7777777777777778
7329.999n 0.3333333333333333 0.6666666666666666 0.0 0.0 0.7777777777777778
7330n 0.3333333333333333 0.0 0.6666666666666666 0.6666666666666666 0.5555555555555556
7339.999n 0.3333333333333333 0.0 0.6666666666666666 0.6666666666666666 0.5555555555555556
7340n 1.0 0.6666666666666666 0.0 1.0 1.4444444444444444
7349.999n 1.0 0.6666666666666666 0.0 1.0 1.4444444444444444
7350n 0.0 0.6666666666666666 1.0 1.0 0.7777777777777778
7359.999n 0.0 0.6666666666666666 1.0 1.0 0.7777777777777778
7360n 0.3333333333333333 1.0 0.0 0.6666666666666666 1.0
7369.999n 0.3333333333333333 1.0 0.0 0.6666666666666666 1.0
7370n 0.6666666666666666 0.6666666666666666 0.3333333333333333 0.6666666666666666 1.2222222222222223
7379.999n 0.6666666666666666 0.6666666666666666 0.3333333333333333 0.6666666666666666 1.2222222222222223
7380n 1.0 0.6666666666666666 0.3333333333333333 0.6666666666666666 1.5555555555555556
7389.999n 1.0 0.6666666666666666 0.3333333333333333 0.6666666666666666 1.5555555555555556
7390n 0.6666666666666666 0.0 0.3333333333333333 0.3333333333333333 0.7777777777777778
7399.999n 0.6666666666666666 0.0 0.3333333333333333 0.3333333333333333 0.7777777777777778
7400n 0.3333333333333333 0.3333333333333333 1.0 0.0 0.8888888888888888
7409.999n 0.3333333333333333 0.3333333333333333 1.0 0.0 0.8888888888888888
7410n 0.0 1.0 0.6666666666666666 0.6666666666666666 0.8888888888888888
7419.999n 0.0 1.0 0.6666666666666666 0.6666666666666666 0.8888888888888888
7420n 0.3333333333333333 0.0 0.6666666666666666 0.3333333333333333 0.5555555555555556
7429.999n 0.3333333333333333 0.0 0.6666666666666666 0.3333333333333333 0.5555555555555556
7430n 0.6666666666666666 0.6666666666666666 1.0 0.6666666666666666 1.4444444444444444
7439.999n 0.6666666666666666 0.6666666666666666 1.0 0.6666666666666666 1.4444444444444444
7440n 0.0 0.6666666666666666 0.6666666666666666 1.0 0.6666666666666666
7449.999n 0.0 0.6666666666666666 0.6666666666666666 1.0 0.6666666666666666
7450n 1.0 0.3333333333333333 0.3333333333333333 1.0 1.3333333333333333
7459.999n 1.0 0.3333333333333333 0.3333333333333333 1.0 1.3333333333333333
7460n 0.3333333333333333 0.0 0.6666666666666666 0.0 0.5555555555555556
7469.999n 0.3333333333333333 0.0 0.6666666666666666 0.0 0.5555555555555556
7470n 0.0 0.0 0.3333333333333333 0.0 0.1111111111111111
7479.999n 0.0 0.0 0.3333333333333333 0.0 0.1111111111111111
7480n 0.6666666666666666 0.6666666666666666 0.0 0.0 1.1111111111111112
7489.999n 0.6666666666666666 0.6666666666666666 0.0 0.0 1.1111111111111112
7490n 0.3333333333333333 1.0 0.0 1.0 1.0
7499.999n 0.3333333333333333 1.0 0.0 1.0 1.0
7500n 1.0 1.0 1.0 0.0 2.0
7509.999n 1.0 1.0 1.0 0.0 2.0
7510n 1.0 1.0 0.6666666666666666 0.6666666666666666 1.8888888888888888
7519.999n 1.0 1.0 0.6666666666666666 0.6666666666666666 1.8888888888888888
7520n 0.0 0.6666666666666666 0.6666666666666666 0.3333333333333333 0.6666666666666666
7529.999n 0.0 0.6666666666666666 0.6666666666666666 0.3333333333333333 0.6666666666666666
7530n 0.0 1.0 0.3333333333333333 0.0 0.7777777777777778
7539.999n 0.0 1.0 0.3333333333333333 0.0 0.7777777777777778
7540n 0.0 0.0 0.6666666666666666 0.0 0.2222222222222222
7549.999n 0.0 0.0 0.6666666666666666 0.0 0.2222222222222222
7550n 0.6666666666666666 1.0 1.0 0.3333333333333333 1.6666666666666667
7559.999n 0.6666666666666666 1.0 1.0 0.3333333333333333 1.6666666666666667
7560n 0.0 1.0 0.0 0.0 0.6666666666666666
7569.999n 0.0 1.0 0.0 0.0 0.6666666666666666
7570n 0.3333333333333333 1.0 0.3333333333333333 0.0 1.1111111111111112
7579.999n 0.3333333333333333 1.0 0.3333333333333333 0.0 1.1111111111111112
7580n 0.3333333333333333 0.3333333333333333 0.3333333333333333 1.0 0.6666666666666666
7589.999n 0.3333333333333333 0.3333333333333333 0.3333333333333333 1.0 0.6666666666666666
7590n 0.0 1.0 1.0 1.0 1.0
7599.999n 0.0 1.0 1.0 1.0 1.0
7600n 1.0 0.6666666666666666 0.6666666666666666 1.0 1.6666666666666667
7609.999n 1.0 0.6666666666666666 0.6666666666666666 1.0 1.6666666666666667
7610n 0.0 0.3333333333333333 0.6666666666666666 0.6666666666666666 0.4444444444444444
7619.999n 0.0 0.3333333333333333 0.6666666666666666 0.6666666666666666 0.4444444444444444
7620n 0.0 1.0 0.6666666666666666 0.0 0.8888888888888888
7629.999n 0.0 1.0 0.6666666666666666 0.0 0.8888888888888888
7630n 0.0 0.0 1.0 1.0 0.3333333333333333
7639.999n 0.0 0.0 1.0 1.0 0.3333333333333333
7640n 0.3333333333333333 0.0 0.3333333333333333 0.6666666666666666 0.4444444444444444
7649.999n 0.3333333333333333 0.0 0.3333333333333333 0.6666666666666666 0.4444444444444444
7650n 0.0 1.0 1.0 0.0 1.0
7659.999n 0.0 1.0 1.0 0.0 1.0
7660n 0.6666666666666666 0.0 1.0 0.3333333333333333 1.0
7669.999n 0.6666666666666666 0.0 1.0 0.3333333333333333 1.0
7670n 0.3333333333333333 0.3333333333333333 0.6666666666666666 0.3333333333333333 0.7777777777777778
7679.999n 0.3333333333333333 0.3333333333333333 0.6666666666666666 0.3333333333333333 0.7777777777777778
7680n 0.3333333333333333 1.0 1.0 0.0 1.3333333333333333
7689.999n 0.3333333333333333 1.0 1.0 0.0 1.3333333333333333
7690n 0.6666666666666666 0.0 0.0 0.6666666666666666 0.6666666666666666
7699.999n 0.6666666666666666 0.0 0.0 0.6666666666666666 0.6666666666666666
7700n 0.6666666666666666 0.6666666666666666 1.0 1.0 1.4444444444444444
7709.999n 0.6666666666666666 0.6666666666666666 1.0 1.0 1.4444444444444444
7710n 0.0 0.0 0.3333333333333333 1.0 0.1111111111111111
7719.999n 0.0 0.0 0.3333333333333333 1.0 0.1111111111111111
7720n 0.3333333333333333 0.6666666666666666 0.6666666666666666 0.6666666666666666 1.0
7729.999n 0.3333333333333333 0.6666666666666666 0.6666666666666666 0.6666666666666666 1.0
7730n 0.3333333333333333 0.6666666666666666 0.3333333333333333 1.0 0.8888888888888888
7739.999n 0.3333333333333333 0.6666666666666666 0.3333333333333333 1.0 0.8888888888888888
7740n 0.3333333333333333 1.0 0.6666666666666666 0.6666666666666666 1.2222222222222223
7749.999n 0.3333333333333333 1.0 0.6666666666666666 0.6666666666666666 1.2222222222222223
7750n 0.0 0.0 0.3333333333333333 1.0 0.1111111111111111
7759.999n 0.0 0.0 0.3333333333333333 1.0 0.1111111111111111
7760n 0.6666666666666666 0.3333333333333333 0.0 0.0 0.8888888888888888
7769.999n 0.6666666666666666 0.3333333333333333 0.0 0.0 0.8888888888888888
7770n 1.0 0.6666666666666666 1.0 0.3333333333333333 1.7777777777777777
7779.999n 1.0 0.6666666666666666 1.0 0.3333333333333333 1.7777777777777777
7780n 1.0 0.3333333333333333 0.6666666666666666 1.0 1.4444444444444444
7789.999n 1.0 0.3333333333333333 0.6666666666666666 1.0 1.4444444444444444
7790n 1.0 0.3333333333333333 0.3333333333333333 0.6666666666666666 1.3333333333333333
7799.999n 1.0 0.3333333333333333 0.3333333333333333 0.6666666666666666 1.3333333333333333
7800n 0.0 0.6666666666666666 0.0 0.6666666666666666 0.4444444444444444
7809.999n 0.0 0.6666666666666666 0.0 0.6666666666666666 0.4444444444444444
7810n 0.0 1.0 0.0 0.6666666666666666 0.6666666666666666
7819.999n 0.0 1.0 0.0 0.6666666666666666 0.6666666666666666
7820n 0.3333333333333333 0.3333333333333333 0.0 0.6666666666666666 0.5555555555555556
7829.999n 0.3333333333333333 0.3333333333333333 0.0 0.6666666666666666 0.5555555555555556
7830n 0.6666666666666666 1.0 0.6666666666666666 0.0 1.5555555555555556
7839.999n 0.6666666666666666 1.0 0.6666666666666666 0.0 1.5555555555555556
7840n 0.6666666666666666 0.3333333333333333 0.3333333333333333 0.3333333333333333 1.0
7849.999n 0.6666666666666666 0.3333333333333333 0.3333333333333333 0.3333333333333333 1.0
7850n 1.0 0.6666666666666666 0.3333333333333333 0.6666666666666666 1.5555555555555556
7859.999n 1.0 0.6666666666666666 0.3333333333333333 0.6666666666666666 1.5555555555555556
7860n 0.3333333333333333 0.0 0.0 0.0 0.3333333333333333
7869.999n 0.3333333333333333 0.0 0.0 0.0 0.3333333333333333
7870n 1.0 0.3333333333333333 0.6666666666666666 1.0 1.4444444444444444
7879.999n 1.0 0.3333333333333333 0.6666666666666666 1.0 1.4444444444444444
7880n 0.6666666666666666 1.0 1.0 0.6666666666666666 1.6666666666666667
7889.999n 0.6666666666666666 1.0 1.0 0.6666666666666666 1.6666666666666667
7890n 0.6666666666666666 0.0 1.0 0.0 1.0
7899.999n 0.6666666666666666 0.0 1.0 0.0 1.0
7900n 1.0 0.0 0.3333333333333333 0.0 1.1111111111111112
7909.999n 1.0 0.0 0.3333333333333333 0.0 1.1111111111111112
7910n 0.3333333333333333 1.0 0.0 0.6666666666666666 1.0
7919.999n 0.3333333333333333 1.0 0.0 0.6666666666666666 1.0
7920n 0.6666666666666666 0.0 0.3333333333333333 0.3333333333333333 0.7777777777777778
7929.999n 0.6666666666666666 0.0 0.3333333333333333 0.3333333333333333 0.7777777777777778
7930n 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.6666666666666666 1.1111111111111112
7939.999n 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.6666666666666666 1.1111111111111112
7940n 0.0 1.0 0.6666666666666666 0.3333333333333333 0.8888888888888888
7949.999n 0.0 1.0 0.6666666666666666 0.3333333333333333 0.8888888888888888
7950n 0.6666666666666666 0.6666666666666666 1.0 0.3333333333333333 1.4444444444444444
7959.999n 0.6666666666666666 0.6666666666666666 1.0 0.3333333333333333 1.4444444444444444
7960n 0.0 0.6666666666666666 0.6666666666666666 0.6666666666666666 0.6666666666666666
7969.999n 0.0 0.6666666666666666 0.6666666666666666 0.6666666666666666 0.6666666666666666
7970n 0.3333333333333333 1.0 1.0 0.0 1.3333333333333333
7979.999n 0.3333333333333333 1.0 1.0 0.0 1.3333333333333333
7980n 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.6666666666666666 1.1111111111111112
7989.999n 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.6666666666666666 1.1111111111111112
7990n 1.0 0.6666666666666666 1.0 1.0 1.7777777777777777
7999.999n 1.0 0.6666666666666666 1.0 1.0 1.7777777777777777
8000n 0.6666666666666666 0.0 0.6666666666666666 0.0 0.8888888888888888
8009.999n 0.6666666666666666 0.0 0.6666666666666666 0.0 0.8888888888888888
8010n 0.6666666666666666 0.0 1.0 0.0 1.0
8019.999n 0.6666666666666666 0.0 1.0 0.0 1.0
8020n 0.0 0.6666666666666666 0.0 0.0 0.4444444444444444
8029.999n 0.0 0.6666666666666666 0.0 0.0 0.4444444444444444
8030n 0.3333333333333333 0.0 1.0 1.0 0.6666666666666666
8039.999n 0.3333333333333333 0.0 1.0 1.0 0.6666666666666666
8040n 0.6666666666666666 1.0 0.3333333333333333 0.6666666666666666 1.4444444444444444
8049.999n 0.6666666666666666 1.0 0.3333333333333333 0.6666666666666666 1.4444444444444444
8050n 0.6666666666666666 1.0 0.3333333333333333 0.6666666666666666 1.4444444444444444
8059.999n 0.6666666666666666 1.0 0.3333333333333333 0.6666666666666666 1.4444444444444444
8060n 0.3333333333333333 0.3333333333333333 0.6666666666666666 0.0 0.7777777777777778
8069.999n 0.3333333333333333 0.3333333333333333 0.6666666666666666 0.0 0.7777777777777778
8070n 0.0 0.3333333333333333 0.0 0.0 0.2222222222222222
8079.999n 0.0 0.3333333333333333 0.0 0.0 0.2222222222222222
8080n 0.0 1.0 0.6666666666666666 0.6666666666666666 0.8888888888888888
8089.999n 0.0 1.0 0.6666666666666666 0.6666666666666666 0.8888888888888888
8090n 0.6666666666666666 0.3333333333333333 0.6666666666666666 1.0 1.1111111111111112
8099.999n 0.6666666666666666 0.3333333333333333 0.6666666666666666 1.0 1.1111111111111112
8100n 1.0 0.3333333333333333 0.0 0.6666666666666666 1.2222222222222223
8109.999n 1.0 0.3333333333333333 0.0 0.6666666666666666 1.2222222222222223
8110n 0.0 0.0 0.0 0.6666666666666666 0.0
8119.999n 0.0 0.0 0.0 0.6666666666666666 0.0
8120n 1.0 1.0 0.6666666666666666 1.0 1.8888888888888888
8129.999n 1.0 1.0 0.6666666666666666 1.0 1.8888888888888888
8130n 1.0 0.0 0.3333333333333333 0.3333333333333333 1.1111111111111112
8139.999n 1.0 0.0 0.3333333333333333 0.3333333333333333 1.1111111111111112
8140n 1.0 0.3333333333333333 0.0 0.0 1.2222222222222223
8149.999n 1.0 0.3333333333333333 0.0 0.0 1.2222222222222223
8150n 1.0 0.0 1.0 0.6666666666666666 1.3333333333333333
8159.999n 1.0 0.0 1.0 0.6666666666666666 1.3333333333333333
8160n 1.0 0.0 0.0 0.0 1.0
8169.999n 1.0 0.0 0.0 0.0 1.0
8170n 0.6666666666666666 0.3333333333333333 0.3333333333333333 0.6666666666666666 1.0
8179.999n 0.6666666666666666 0.3333333333333333 0.3333333333333333 0.6666666666666666 1.0
8180n 1.0 1.0 0.6666666666666666 0.6666666666666666 1.8888888888888888
8189.999n 1.0 1.0 0.6666666666666666 0.6666666666666666 1.8888888888888888
8190n 0.3333333333333333 0.3333333333333333 1.0 0.0 0.8888888888888888
8199.999n 0.3333333333333333 0.3333333333333333 1.0 0.0 0.8888888888888888
8200n 1.0 0.6666666666666666 0.6666666666666666 0.0 1.6666666666666667
8209.999n 1.0 0.6666666666666666 0.6666666666666666 0.0 1.6666666666666667
8210n 0.3333333333333333 0.0 1.0 0.0 0.6666666666666666
8219.999n 0.3333333333333333 0.0 1.0 0.0 0.6666666666666666
8220n 1.0 1.0 0.0 0.0 1.6666666666666667
8229.999n 1.0 1.0 0.0 0.0 1.6666666666666667
8230n 0.3333333333333333 1.0 1.0 0.6666666666666666 1.3333333333333333
8239.999n 0.3333333333333333 1.0 1.0 0.6666666666666666 1.3333333333333333
8240n 0.6666666666666666 1.0 1.0 1.0 1.6666666666666667
8249.999n 0.6666666666666666 1.0 1.0 1.0 1.6666666666666667
8250n 0.3333333333333333 0.6666666666666666 0.6666666666666666 0.3333333333333333 1.0
8259.999n 0.3333333333333333 0.6666666666666666 0.6666666666666666 0.3333333333333333 1.0
8260n 1.0 0.6666666666666666 0.0 0.0 1.4444444444444444
8269.999n 1.0 0.6666666666666666 0.0 0.0 1.4444444444444444
8270n 0.6666666666666666 1.0 0.3333333333333333 0.0 1.4444444444444444
8279.999n 0.6666666666666666 1.0 0.3333333333333333 0.0 1.4444444444444444
8280n 0.6666666666666666 1.0 0.3333333333333333 0.3333333333333333 1.4444444444444444
8289.999n 0.6666666666666666 1.0 0.3333333333333333 0.3333333333333333 1.4444444444444444
8290n 0.3333333333333333 0.6666666666666666 0.6666666666666666 0.6666666666666666 1.0
8299.999n 0.3333333333333333 0.6666666666666666 0.6666666666666666 0.6666666666666666 1.0
8300n 1.0 0.3333333333333333 0.0 1.0 1.2222222222222223
8309.999n 1.0 0.3333333333333333 0.0 1.0 1.2222222222222223
8310n 0.3333333333333333 0.0 1.0 0.0 0.6666666666666666
8319.999n 0.3333333333333333 0.0 1.0 0.0 0.6666666666666666
8320n 0.3333333333333333 1.0 1.0 1.0 1.3333333333333333
8329.999n 0.3333333333333333 1.0 1.0 1.0 1.3333333333333333
8330n 1.0 1.0 0.0 0.0 1.6666666666666667
8339.999n 1.0 1.0 0.0 0.0 1.6666666666666667
8340n 0.3333333333333333 0.0 0.6666666666666666 0.0 0.5555555555555556
8349.999n 0.3333333333333333 0.0 0.6666666666666666 0.0 0.5555555555555556
8350n 0.0 0.0 1.0 0.3333333333333333 0.3333333333333333
8359.999n 0.0 0.0 1.0 0.3333333333333333 0.3333333333333333
8360n 0.0 0.3333333333333333 0.0 0.3333333333333333 0.2222222222222222
8369.999n 0.0 0.3333333333333333 0.0 0.3333333333333333 0.2222222222222222
8370n 0.6666666666666666 1.0 0.3333333333333333 0.0 1.4444444444444444
8379.999n 0.6666666666666666 1.0 0.3333333333333333 0.0 1.4444444444444444
8380n 0.0 1.0 0.3333333333333333 0.3333333333333333 0.7777777777777778
8389.999n 0.0 1.0 0.3333333333333333 0.3333333333333333 0.7777777777777778
8390n 0.3333333333333333 0.3333333333333333 0.6666666666666666 0.0 0.7777777777777778
8399.999n 0.3333333333333333 0.3333333333333333 0.6666666666666666 0.0 0.7777777777777778
8400n 0.6666666666666666 1.0 0.3333333333333333 0.6666666666666666 1.4444444444444444
8409.999n 0.6666666666666666 1.0 0.3333333333333333 0.6666666666666666 1.4444444444444444
8410n 0.0 0.3333333333333333 0.3333333333333333 0.0 0.3333333333333333
8419.999n 0.0 0.3333333333333333 0.3333333333333333 0.0 0.3333333333333333
8420n 0.0 1.0 1.0 1.0 1.0
8429.999n 0.0 1.0 1.0 1.0 1.0
8430n 1.0 1.0 1.0 1.0 2.0
8439.999n 1.0 1.0 1.0 1.0 2.0
8440n 0.0 1.0 0.3333333333333333 1.0 0.7777777777777778
8449.999n 0.0 1.0 0.3333333333333333 1.0 0.7777777777777778
8450n 1.0 0.3333333333333333 1.0 1.0 1.5555555555555556
8459.999n 1.0 0.3333333333333333 1.0 1.0 1.5555555555555556
8460n 1.0 0.3333333333333333 1.0 0.6666666666666666 1.5555555555555556
8469.999n 1.0 0.3333333333333333 1.0 0.6666666666666666 1.5555555555555556
8470n 1.0 1.0 0.6666666666666666 0.3333333333333333 1.8888888888888888
8479.999n 1.0 1.0 0.6666666666666666 0.3333333333333333 1.8888888888888888
8480n 0.0 1.0 1.0 0.6666666666666666 1.0
8489.999n 0.0 1.0 1.0 0.6666666666666666 1.0
8490n 0.6666666666666666 0.3333333333333333 1.0 0.3333333333333333 1.2222222222222223
8499.999n 0.6666666666666666 0.3333333333333333 1.0 0.3333333333333333 1.2222222222222223
8500n 0.0 0.0 0.6666666666666666 0.6666666666666666 0.2222222222222222
8509.999n 0.0 0.0 0.6666666666666666 0.6666666666666666 0.2222222222222222
8510n 1.0 1.0 0.0 0.3333333333333333 1.6666666666666667
8519.999n 1.0 1.0 0.0 0.3333333333333333 1.6666666666666667
8520n 0.3333333333333333 1.0 1.0 0.0 1.3333333333333333
8529.999n 0.3333333333333333 1.0 1.0 0.0 1.3333333333333333
8530n 0.3333333333333333 0.3333333333333333 1.0 0.0 0.8888888888888888
8539.999n 0.3333333333333333 0.3333333333333333 1.0 0.0 0.8888888888888888
8540n 0.3333333333333333 0.6666666666666666 0.0 1.0 0.7777777777777778
8549.999n 0.3333333333333333 0.6666666666666666 0.0 1.0 0.7777777777777778
8550n 0.3333333333333333 0.3333333333333333 0.0 1.0 0.5555555555555556
8559.999n 0.3333333333333333 0.3333333333333333 0.0 1.0 0.5555555555555556
8560n 0.3333333333333333 1.0 0.3333333333333333 0.3333333333333333 1.1111111111111112
8569.999n 0.3333333333333333 1.0 0.3333333333333333 0.3333333333333333 1.1111111111111112
8570n 0.0 1.0 0.6666666666666666 1.0 0.8888888888888888
8579.999n 0.0 1.0 0.6666666666666666 1.0 0.8888888888888888
8580n 1.0 1.0 0.6666666666666666 1.0 1.8888888888888888
8589.999n 1.0 1.0 0.6666666666666666 1.0 1.8888888888888888
8590n 0.3333333333333333 0.6666666666666666 0.6666666666666666 1.0 1.0
8599.999n 0.3333333333333333 0.6666666666666666 0.6666666666666666 1.0 1.0
8600n 0.0 0.3333333333333333 1.0 0.3333333333333333 0.5555555555555556
8609.999n 0.0 0.3333333333333333 1.0 0.3333333333333333 0.5555555555555556
8610n 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.6666666666666666 1.1111111111111112
8619.999n 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.6666666666666666 1.1111111111111112
8620n 0.0 1.0 0.6666666666666666 0.3333333333333333 0.8888888888888888
8629.999n 0.0 1.0 0.6666666666666666 0.3333333333333333 0.8888888888888888
8630n 0.6666666666666666 0.6666666666666666 0.6666666666666666 1.0 1.3333333333333333
8639.999n 0.6666666666666666 0.6666666666666666 0.6666666666666666 1.0 1.3333333333333333
8640n 0.3333333333333333 0.3333333333333333 0.3333333333333333 1.0 0.6666666666666666
8649.999n 0.3333333333333333 0.3333333333333333 0.3333333333333333 1.0 0.6666666666666666
8650n 1.0 0.3333333333333333 0.6666666666666666 1.0 1.4444444444444444
8659.999n 1.0 0.3333333333333333 0.6666666666666666 1.0 1.4444444444444444
8660n 1.0 1.0 0.3333333333333333 0.3333333333333333 1.7777777777777777
8669.999n 1.0 1.0 0.3333333333333333 0.3333333333333333 1.7777777777777777
8670n 0.0 0.0 1.0 0.6666666666666666 0.3333333333333333
8679.999n 0.0 0.0 1.0 0.6666666666666666 0.3333333333333333
8680n 0.0 1.0 0.0 1.0 0.6666666666666666
8689.999n 0.0 1.0 0.0 1.0 0.6666666666666666
8690n 1.0 0.6666666666666666 0.3333333333333333 0.0 1.5555555555555556
8699.999n 1.0 0.6666666666666666 0.3333333333333333 0.0 1.5555555555555556
8700n 0.3333333333333333 1.0 1.0 0.0 1.3333333333333333
8709.999n 0.3333333333333333 1.0 1.0 0.0 1.3333333333333333
8710n 0.3333333333333333 0.6666666666666666 0.6666666666666666 0.3333333333333333 1.0
8719.999n 0.3333333333333333 0.6666666666666666 0.6666666666666666 0.3333333333333333 1.0
8720n 0.6666666666666666 0.3333333333333333 0.0 0.0 0.8888888888888888
8729.999n 0.6666666666666666 0.3333333333333333 0.0 0.0 0.8888888888888888
8730n 0.6666666666666666 0.0 0.0 1.0 0.6666666666666666
8739.999n 0.6666666666666666 0.0 0.0 1.0 0.6666666666666666
8740n 0.6666666666666666 1.0 1.0 0.0 1.6666666666666667
8749.999n 0.6666666666666666 1.0 1.0 0.0 1.6666666666666667
8750n 0.6666666666666666 0.6666666666666666 0.6666666666666666 1.0 1.3333333333333333
8759.999n 0.6666666666666666 0.6666666666666666 0.6666666666666666 1.0 1.3333333333333333
8760n 0.6666666666666666 0.0 0.0 0.0 0.6666666666666666
8769.999n 0.6666666666666666 0.0 0.0 0.0 0.6666666666666666
8770n 0.0 0.0 0.3333333333333333 0.0 0.1111111111111111
8779.999n 0.0 0.0 0.3333333333333333 0.0 0.1111111111111111
8780n 0.6666666666666666 0.6666666666666666 0.0 0.3333333333333333 1.1111111111111112
8789.999n 0.6666666666666666 0.6666666666666666 0.0 0.3333333333333333 1.1111111111111112
8790n 1.0 1.0 1.0 0.0 2.0
8799.999n 1.0 1.0 1.0 0.0 2.0
8800n 0.3333333333333333 1.0 0.3333333333333333 0.6666666666666666 1.1111111111111112
8809.999n 0.3333333333333333 1.0 0.3333333333333333 0.6666666666666666 1.1111111111111112
8810n 1.0 0.6666666666666666 0.3333333333333333 0.0 1.5555555555555556
8819.999n 1.0 0.6666666666666666 0.3333333333333333 0.0 1.5555555555555556
8820n 0.3333333333333333 1.0 0.3333333333333333 0.0 1.1111111111111112
8829.999n 0.3333333333333333 1.0 0.3333333333333333 0.0 1.1111111111111112
8830n 0.6666666666666666 0.6666666666666666 0.3333333333333333 0.0 1.2222222222222223
8839.999n 0.6666666666666666 0.6666666666666666 0.3333333333333333 0.0 1.2222222222222223
8840n 0.6666666666666666 1.0 0.6666666666666666 0.0 1.5555555555555556
8849.999n 0.6666666666666666 1.0 0.6666666666666666 0.0 1.5555555555555556
8850n 0.0 0.3333333333333333 0.0 0.3333333333333333 0.2222222222222222
8859.999n 0.0 0.3333333333333333 0.0 0.3333333333333333 0.2222222222222222
8860n 0.0 0.0 0.0 0.3333333333333333 0.0
8869.999n 0.0 0.0 0.0 0.3333333333333333 0.0
8870n 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.6666666666666666 1.1111111111111112
8879.999n 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.6666666666666666 1.1111111111111112
8880n 0.3333333333333333 1.0 1.0 0.3333333333333333 1.3333333333333333
8889.999n 0.3333333333333333 1.0 1.0 0.3333333333333333 1.3333333333333333
8890n 0.3333333333333333 0.0 0.3333333333333333 0.3333333333333333 0.4444444444444444
8899.999n 0.3333333333333333 0.0 0.3333333333333333 0.3333333333333333 0.4444444444444444
8900n 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.0 1.1111111111111112
8909.999n 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.0 1.1111111111111112
8910n 0.3333333333333333 0.0 1.0 0.6666666666666666 0.6666666666666666
8919.999n 0.3333333333333333 0.0 1.0 0.6666666666666666 0.6666666666666666
8920n 0.6666666666666666 0.0 0.3333333333333333 0.0 0.7777777777777778
8929.999n 0.6666666666666666 0.0 0.3333333333333333 0.0 0.7777777777777778
8930n 0.3333333333333333 1.0 0.3333333333333333 0.0 1.1111111111111112
8939.999n 0.3333333333333333 1.0 0.3333333333333333 0.0 1.1111111111111112
8940n 1.0 0.6666666666666666 0.6666666666666666 0.6666666666666666 1.6666666666666667
8949.999n 1.0 0.6666666666666666 0.6666666666666666 0.6666666666666666 1.6666666666666667
8950n 1.0 0.6666666666666666 0.0 1.0 1.4444444444444444
8959.999n 1.0 0.6666666666666666 0.0 1.0 1.4444444444444444
8960n 0.6666666666666666 0.6666666666666666 0.0 1.0 1.1111111111111112
8969.999n 0.6666666666666666 0.6666666666666666 0.0 1.0 1.1111111111111112
8970n 0.3333333333333333 0.6666666666666666 0.3333333333333333 0.0 0.8888888888888888
8979.999n 0.3333333333333333 0.6666666666666666 0.3333333333333333 0.0 0.8888888888888888
8980n 0.0 0.3333333333333333 0.3333333333333333 0.6666666666666666 0.3333333333333333
8989.999n 0.0 0.3333333333333333 0.3333333333333333 0.6666666666666666 0.3333333333333333
8990n 0.6666666666666666 0.3333333333333333 0.0 0.0 0.8888888888888888
8999.999n 0.6666666666666666 0.3333333333333333 0.0 0.0 0.8888888888888888
9000n 0.6666666666666666 1.0 0.6666666666666666 0.3333333333333333 1.5555555555555556
9009.999n 0.6666666666666666 1.0 0.6666666666666666 0.3333333333333333 1.5555555555555556
9010n 0.3333333333333333 0.3333333333333333 0.6666666666666666 0.3333333333333333 0.7777777777777778
9019.999n 0.3333333333333333 0.3333333333333333 0.6666666666666666 0.3333333333333333 0.7777777777777778
9020n 1.0 0.0 0.3333333333333333 0.3333333333333333 1.1111111111111112
9029.999n 1.0 0.0 0.3333333333333333 0.3333333333333333 1.1111111111111112
9030n 0.0 0.6666666666666666 1.0 0.3333333333333333 0.7777777777777778
9039.999n 0.0 0.6666666666666666 1.0 0.3333333333333333 0.7777777777777778
9040n 1.0 1.0 0.6666666666666666 0.3333333333333333 1.8888888888888888
9049.999n 1.0 1.0 0.6666666666666666 0.3333333333333333 1.8888888888888888
9050n 0.0 0.3333333333333333 0.3333333333333333 1.0 0.3333333333333333
9059.999n 0.0 0.3333333333333333 0.3333333333333333 1.0 0.3333333333333333
9060n 0.6666666666666666 0.6666666666666666 0.3333333333333333 0.6666666666666666 1.2222222222222223
9069.999n 0.6666666666666666 0.6666666666666666 0.3333333333333333 0.6666666666666666 1.2222222222222223
9070n 0.0 0.6666666666666666 0.0 1.0 0.4444444444444444
9079.999n 0.0 0.6666666666666666 0.0 1.0 0.4444444444444444
9080n 1.0 0.3333333333333333 0.6666666666666666 1.0 1.4444444444444444
9089.999n 1.0 0.3333333333333333 0.6666666666666666 1.0 1.4444444444444444
9090n 0.6666666666666666 1.0 1.0 0.6666666666666666 1.6666666666666667
9099.999n 0.6666666666666666 1.0 1.0 0.6666666666666666 1.6666666666666667
9100n 0.3333333333333333 1.0 0.0 0.6666666666666666 1.0
9109.999n 0.3333333333333333 1.0 0.0 0.6666666666666666 1.0
9110n 0.6666666666666666 0.6666666666666666 1.0 0.0 1.4444444444444444
9119.999n 0.6666666666666666 0.6666666666666666 1.0 0.0 1.4444444444444444
9120n 1.0 0.0 0.3333333333333333 1.0 1.1111111111111112
9129.999n 1.0 0.0 0.3333333333333333 1.0 1.1111111111111112
9130n 0.6666666666666666 1.0 0.0 1.0 1.3333333333333333
9139.999n 0.6666666666666666 1.0 0.0 1.0 1.3333333333333333
9140n 0.0 0.6666666666666666 0.0 0.6666666666666666 0.4444444444444444
9149.999n 0.0 0.6666666666666666 0.0 0.6666666666666666 0.4444444444444444
9150n 1.0 0.6666666666666666 1.0 0.0 1.7777777777777777
9159.999n 1.0 0.6666666666666666 1.0 0.0 1.7777777777777777
9160n 0.0 0.3333333333333333 0.0 1.0 0.2222222222222222
9169.999n 0.0 0.3333333333333333 0.0 1.0 0.2222222222222222
9170n 0.6666666666666666 0.3333333333333333 1.0 0.6666666666666666 1.2222222222222223
9179.999n 0.6666666666666666 0.3333333333333333 1.0 0.6666666666666666 1.2222222222222223
9180n 0.6666666666666666 0.3333333333333333 0.0 1.0 0.8888888888888888
9189.999n 0.6666666666666666 0.3333333333333333 0.0 1.0 0.8888888888888888
9190n 0.3333333333333333 0.6666666666666666 0.0 0.0 0.7777777777777778
9199.999n 0.3333333333333333 0.6666666666666666 0.0 0.0 0.7777777777777778
9200n 0.3333333333333333 1.0 0.6666666666666666 0.6666666666666666 1.2222222222222223
9209.999n 0.3333333333333333 1.0 0.6666666666666666 0.6666666666666666 1.2222222222222223
9210n 0.6666666666666666 0.6666666666666666 0.3333333333333333 0.3333333333333333 1.2222222222222223
9219.999n 0.6666666666666666 0.6666666666666666 0.3333333333333333 0.3333333333333333 1.2222222222222223
9220n 0.0 0.3333333333333333 0.6666666666666666 0.0 0.4444444444444444
9229.999n 0.0 0.3333333333333333 0.6666666666666666 0.0 0.4444444444444444
9230n 1.0 0.0 0.3333333333333333 0.3333333333333333 1.1111111111111112
9239.999n 1.0 0.0 0.3333333333333333 0.3333333333333333 1.1111111111111112
9240n 0.6666666666666666 0.0 1.0 0.6666666666666666 1.0
9249.999n 0.6666666666666666 0.0 1.0 0.6666666666666666 1.0
9250n 0.6666666666666666 0.3333333333333333 0.6666666666666666 1.0 1.1111111111111112
9259.999n 0.6666666666666666 0.3333333333333333 0.6666666666666666 1.0 1.1111111111111112
9260n 0.6666666666666666 0.0 1.0 0.0 1.0
9269.999n 0.6666666666666666 0.0 1.0 0.0 1.0
9270n 0.6666666666666666 0.3333333333333333 1.0 1.0 1.2222222222222223
9279.999n 0.6666666666666666 0.3333333333333333 1.0 1.0 1.2222222222222223
9280n 0.3333333333333333 0.6666666666666666 0.6666666666666666 0.6666666666666666 1.0
9289.999n 0.3333333333333333 0.6666666666666666 0.6666666666666666 0.6666666666666666 1.0
9290n 0.0 0.3333333333333333 0.3333333333333333 0.6666666666666666 0.3333333333333333
9299.999n 0.0 0.3333333333333333 0.3333333333333333 0.6666666666666666 0.3333333333333333
9300n 0.3333333333333333 0.3333333333333333 0.6666666666666666 0.3333333333333333 0.7777777777777778
9309.999n 0.3333333333333333 0.3333333333333333 0.6666666666666666 0.3333333333333333 0.7777777777777778
9310n 0.6666666666666666 0.0 0.6666666666666666 1.0 0.8888888888888888
9319.999n 0.6666666666666666 0.0 0.6666666666666666 1.0 0.8888888888888888
9320n 1.0 0.6666666666666666 0.3333333333333333 1.0 1.5555555555555556
9329.999n 1.0 0.6666666666666666 0.3333333333333333 1.0 1.5555555555555556
9330n 0.0 0.6666666666666666 0.3333333333333333 1.0 0.5555555555555556
9339.999n 0.0 0.6666666666666666 0.3333333333333333 1.0 0.5555555555555556
9340n 0.0 0.6666666666666666 0.3333333333333333 0.3333333333333333 0.5555555555555556
9349.999n 0.0 0.6666666666666666 0.3333333333333333 0.3333333333333333 0.5555555555555556
9350n 1.0 0.3333333333333333 0.6666666666666666 0.3333333333333333 1.4444444444444444
9359.999n 1.0 0.3333333333333333 0.6666666666666666 0.3333333333333333 1.4444444444444444
9360n 0.3333333333333333 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.8888888888888888
9369.999n 0.3333333333333333 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.8888888888888888
9370n 0.0 0.6666666666666666 0.3333333333333333 0.3333333333333333 0.5555555555555556
9379.999n 0.0 0.6666666666666666 0.3333333333333333 0.3333333333333333 0.5555555555555556
9380n 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.6666666666666666 1.1111111111111112
9389.999n 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.6666666666666666 1.1111111111111112
9390n 0.0 0.6666666666666666 0.3333333333333333 1.0 0.5555555555555556
9399.999n 0.0 0.6666666666666666 0.3333333333333333 1.0 0.5555555555555556
9400n 0.6666666666666666 1.0 0.6666666666666666 0.3333333333333333 1.5555555555555556
9409.999n 0.6666666666666666 1.0 0.6666666666666666 0.3333333333333333 1.5555555555555556
9410n 0.3333333333333333 0.0 1.0 1.0 0.6666666666666666
9419.999n 0.3333333333333333 0.0 1.0 1.0 0.6666666666666666
9420n 1.0 1.0 1.0 0.0 2.0
9429.999n 1.0 1.0 1.0 0.0 2.0
9430n 0.3333333333333333 0.0 0.0 0.3333333333333333 0.3333333333333333
9439.999n 0.3333333333333333 0.0 0.0 0.3333333333333333 0.3333333333333333
9440n 0.0 0.6666666666666666 0.0 0.6666666666666666 0.4444444444444444
9449.999n 0.0 0.6666666666666666 0.0 0.6666666666666666 0.4444444444444444
9450n 0.0 0.3333333333333333 1.0 0.3333333333333333 0.5555555555555556
9459.999n 0.0 0.3333333333333333 1.0 0.3333333333333333 0.5555555555555556
9460n 0.0 1.0 0.3333333333333333 0.6666666666666666 0.7777777777777778
9469.999n 0.0 1.0 0.3333333333333333 0.6666666666666666 0.7777777777777778
9470n 0.3333333333333333 0.6666666666666666 1.0 1.0 1.1111111111111112
9479.999n 0.3333333333333333 0.6666666666666666 1.0 1.0 1.1111111111111112
9480n 0.6666666666666666 0.0 0.3333333333333333 0.3333333333333333 0.7777777777777778
9489.999n 0.6666666666666666 0.0 0.3333333333333333 0.3333333333333333 0.7777777777777778
9490n 0.3333333333333333 0.6666666666666666 0.6666666666666666 0.6666666666666666 1.0
9499.999n 0.3333333333333333 0.6666666666666666 0.6666666666666666 0.6666666666666666 1.0
9500n 1.0 1.0 1.0 1.0 2.0
9509.999n 1.0 1.0 1.0 1.0 2.0
9510n 0.6666666666666666 1.0 0.3333333333333333 0.6666666666666666 1.4444444444444444
9519.999n 0.6666666666666666 1.0 0.3333333333333333 0.6666666666666666 1.4444444444444444
9520n 0.3333333333333333 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.8888888888888888
9529.999n 0.3333333333333333 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.8888888888888888
9530n 0.3333333333333333 0.6666666666666666 0.6666666666666666 0.0 1.0
9539.999n 0.3333333333333333 0.6666666666666666 0.6666666666666666 0.0 1.0
9540n 0.6666666666666666 1.0 1.0 0.0 1.6666666666666667
9549.999n 0.6666666666666666 1.0 1.0 0.0 1.6666666666666667
9550n 0.3333333333333333 0.0 1.0 1.0 0.6666666666666666
9559.999n 0.3333333333333333 0.0 1.0 1.0 0.6666666666666666
9560n 0.0 0.3333333333333333 1.0 0.3333333333333333 0.5555555555555556
9569.999n 0.0 0.3333333333333333 1.0 0.3333333333333333 0.5555555555555556
9570n 0.6666666666666666 0.0 1.0 0.0 1.0
9579.999n 0.6666666666666666 0.0 1.0 0.0 1.0
9580n 1.0 0.0 1.0 0.3333333333333333 1.3333333333333333
9589.999n 1.0 0.0 1.0 0.3333333333333333 1.3333333333333333
9590n 0.3333333333333333 0.0 0.0 0.0 0.3333333333333333
9599.999n 0.3333333333333333 0.0 0.0 0.0 0.3333333333333333
9600n 1.0 0.3333333333333333 0.3333333333333333 0.6666666666666666 1.3333333333333333
9609.999n 1.0 0.3333333333333333 0.3333333333333333 0.6666666666666666 1.3333333333333333
9610n 1.0 0.6666666666666666 1.0 0.6666666666666666 1.7777777777777777
9619.999n 1.0 0.6666666666666666 1.0 0.6666666666666666 1.7777777777777777
9620n 0.6666666666666666 0.6666666666666666 1.0 0.3333333333333333 1.4444444444444444
9629.999n 0.6666666666666666 0.6666666666666666 1.0 0.3333333333333333 1.4444444444444444
9630n 0.6666666666666666 1.0 0.3333333333333333 1.0 1.4444444444444444
9639.999n 0.6666666666666666 1.0 0.3333333333333333 1.0 1.4444444444444444
9640n 0.0 0.0 0.3333333333333333 0.3333333333333333 0.1111111111111111
9649.999n 0.0 0.0 0.3333333333333333 0.3333333333333333 0.1111111111111111
9650n 0.3333333333333333 0.3333333333333333 0.3333333333333333 0.3333333333333333 0.6666666666666666
9659.999n 0.3333333333333333 0.3333333333333333 0.3333333333333333 0.3333333333333333 0.6666666666666666
9660n 0.6666666666666666 1.0 0.6666666666666666 0.3333333333333333 1.5555555555555556
9669.999n 0.6666666666666666 1.0 0.6666666666666666 0.3333333333333333 1.5555555555555556
9670n 0.6666666666666666 0.6666666666666666 0.6666666666666666 0.6666666666666666 1.3333333333333333
9679.999n 0.6666666666666666 0.6666666666666666 0.6666666666666666 0.6666666666666666 1.3333333333333333
9680n 0.3333333333333333 0.3333333333333333 0.0 1.0 0.5555555555555556
9689.999n 0.3333333333333333 0.3333333333333333 0.0 1.0 0.5555555555555556
9690n 0.0 1.0 0.6666666666666666 0.6666666666666666 0.8888888888888888
9699.999n 0.0 1.0 0.6666666666666666 0.6666666666666666 0.8888888888888888
9700n 0.3333333333333333 0.3333333333333333 0.6666666666666666 0.3333333333333333 0.7777777777777778
9709.999n 0.3333333333333333 0.3333333333333333 0.6666666666666666 0.3333333333333333 0.7777777777777778
9710n 0.0 0.6666666666666666 0.6666666666666666 1.0 0.6666666666666666
9719.999n 0.0 0.6666666666666666 0.6666666666666666 1.0 0.6666666666666666
9720n 0.0 1.0 1.0 0.3333333333333333 1.0
9729.999n 0.0 1.0 1.0 0.3333333333333333 1.0
9730n 0.3333333333333333 1.0 1.0 0.6666666666666666 1.3333333333333333
9739.999n 0.3333333333333333 1.0 1.0 0.6666666666666666 1.3333333333333333
9740n 0.6666666666666666 0.0 0.3333333333333333 1.0 0.7777777777777778
9749.999n 0.6666666666666666 0.0 0.3333333333333333 1.0 0.7777777777777778
9750n 0.6666666666666666 0.0 0.3333333333333333 0.0 0.7777777777777778
9759.999n 0.6666666666666666 0.0 0.3333333333333333 0.0 0.7777777777777778
9760n 0.3333333333333333 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.8888888888888888
9769.999n 0.3333333333333333 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.8888888888888888
9770n 1.0 0.0 0.6666666666666666 0.3333333333333333 1.2222222222222223
9779.999n 1.0 0.0 0.6666666666666666 0.3333333333333333 1.2222222222222223
9780n 1.0 0.6666666666666666 0.6666666666666666 0.0 1.6666666666666667
9789.999n 1.0 0.6666666666666666 0.6666666666666666 0.0 1.6666666666666667
9790n 1.0 0.6666666666666666 0.3333333333333333 1.0 1.5555555555555556
9799.999n 1.0 0.6666666666666666 0.3333333333333333 1.0 1.5555555555555556
9800n 0.0 0.0 0.3333333333333333 0.6666666666666666 0.1111111111111111
9809.999n 0.0 0.0 0.3333333333333333 0.6666666666666666 0.1111111111111111
9810n 1.0 0.6666666666666666 1.0 0.0 1.7777777777777777
9819.999n 1.0 0.6666666666666666 1.0 0.0 1.7777777777777777
9820n 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.3333333333333333 1.1111111111111112
9829.999n 0.6666666666666666 0.3333333333333333 0.6666666666666666 0.3333333333333333 1.1111111111111112
9830n 0.6666666666666666 0.6666666666666666 0.6666666666666666 0.6666666666666666 1.3333333333333333
9839.999n 0.6666666666666666 0.6666666666666666 0.6666666666666666 0.6666666666666666 1.3333333333333333
9840n 1.0 1.0 0.6666666666666666 0.6666666666666666 1.8888888888888888
9849.999n 1.0 1.0 0.6666666666666666 0.6666666666666666 1.8888888888888888
9850n 0.0 0.0 0.0 1.0 0.0
9859.999n 0.0 0.0 0.0 1.0 0.0
9860n 1.0 0.6666666666666666 0.3333333333333333 0.3333333333333333 1.5555555555555556
9869.999n 1.0 0.6666666666666666 0.3333333333333333 0.3333333333333333 1.5555555555555556
9870n 0.0 1.0 0.0 0.6666666666666666 0.6666666666666666
9879.999n 0.0 1.0 0.0 0.6666666666666666 0.6666666666666666
9880n 0.6666666666666666 0.6666666666666666 0.3333333333333333 1.0 1.2222222222222223
9889.999n 0.6666666666666666 0.6666666666666666 0.3333333333333333 1.0 1.2222222222222223
9890n 0.6666666666666666 0.0 0.0 0.0 0.6666666666666666
9899.999n 0.6666666666666666 0.0 0.0 0.0 0.6666666666666666
9900n 0.3333333333333333 0.0 0.6666666666666666 0.6666666666666666 0.5555555555555556
9909.999n 0.3333333333333333 0.0 0.6666666666666666 0.6666666666666666 0.5555555555555556
9910n 1.0 0.6666666666666666 1.0 1.0 1.7777777777777777
9919.999n 1.0 0.6666666666666666 1.0 1.0 1.7777777777777777
9920n 1.0 0.6666666666666666 0.0 0.6666666666666666 1.4444444444444444
9929.999n 1.0 0.6666666666666666 0.0 0.6666666666666666 1.4444444444444444
9930n 0.0 0.0 1.0 0.3333333333333333 0.3333333333333333
9939.999n 0.0 0.0 1.0 0.3333333333333333 0.3333333333333333
9940n 0.0 0.6666666666666666 0.0 0.0 0.4444444444444444
9949.999n 0.0 0.6666666666666666 0.0 0.0 0.4444444444444444
9950n 0.3333333333333333 0.3333333333333333 0.6666666666666666 0.0 0.7777777777777778
9959.999n 0.3333333333333333 0.3333333333333333 0.6666666666666666 0.0 0.7777777777777778
9960n 1.0 1.0 0.3333333333333333 0.6666666666666666 1.7777777777777777
9969.999n 1.0 1.0 0.3333333333333333 0.6666666666666666 1.7777777777777777
9970n 0.3333333333333333 0.0 0.0 0.3333333333333333 0.3333333333333333
9979.999n 0.3333333333333333 0.0 0.0 0.3333333333333333 0.3333333333333333
9980n 0.6666666666666666 0.6666666666666666 0.0 0.6666666666666666 1.1111111111111112
9989.999n 0.6666666666666666 0.6666666666666666 0.0 0.6666666666666666 1.1111111111111112
9990n 0.3333333333333333 0.0 0.0 0.6666666666666666 0.3333333333333333
9999.999n 0.3333333333333333 0.0 0.0 0.6666666666666666 0.3333333333333333
10000n 0 0 0 0 0
10009.999n 0 0 0 0 0
10010n 1 1 1 1 2
10019.999n 1 1 1 1 2
10020n 0 0 0 0 0
10030n 0 0 0 0 0
.ENDDATA
.TRAN DATA=vector

.measure tran avgpower            AVG power            from=0n to=10030n
.measure tran avg_error           AVG V(expected,Vo) from=0n to=10030n
.measure tran avg_expected_output AVG V(expected)      from=0n to=10030n
.measure tran t0000_1111 trig V(BL1) td=10005n val=0.5 cross=1 targ V(Vo) td=10005n val=1 cross=1
.measure tran t1111_0000 trig V(BL1) td=10015n val=0.5 cross=1 targ V(Vo) td=10015n val=1 cross=1

V_SL1_SET    SL1   0   PWL   0n 0
V_SLref      SLref 0   PWL   0n 0
V_WL         WL    0   PWL   0n 1

.plot tran V(expected, Vo)
.plot tran error = par('V(expected, Vo)/V(expected)*100')
.end